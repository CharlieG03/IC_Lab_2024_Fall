`define CYCLE_TIME 10 // Cycle time in nanoseconds
`define PAT_NUM 10000    // Number of patterns

module PATTERN
`protected
]b3a,ID=Qea4B6;a]eGgFfI5.4)XQ#B1b24;U[NUSOT;(:0K+7JO))&6N]gTT\d5
WfB#Q9O43dUH=.8+]D-==QCM3ISa0OUOB>WO]:1GE^EB/(8=0O4WDK_/<HgA6TgR
>EU^TR&7K9XJG(Y0PU3(>(/#H5T<\W0QL&-.GPg@48S\2,JW)Wd/4b#.;YdAEcbR
KXR^JNb40VXa&fg=+Q\6#F,4M@gQ3Ne7MeEV\9CZK0aQ&RGQ8JbEL:.fX1]1WUQ9
-c>;YK(+1e?3HQ3F-+,X^E/WQR7<E]G/7XEY<H]N>^ZK)c<A.#@4>4=K8Jd[9C]&
?#eYCf_ef1F,P=GgA?1U?M@\/#)D]9BR(ABENE0Y<c6>dcG&fBU&\)[cQgE@:UM.
_Q>OLZBfRRV;E2Ad^2L8O/E;A8Z.]>4a\<U0\UEF@K+CC7=Y137((?;H<8K@#/f>
6A<RQ6@@]fVY70Q2E?F@7819?0Z^>SF5(F=Q0IRI@5#EUJfg/NI,FQ;E-992@&+9
A5Kd8=);1A04UeU)D#D:fNGS7gL]B:_&D,W/>dL;,U2G/RM7TL6>fCgZd3CJNVYg
[OXS;]/(==><H,81O7N@dHC[6Y?D)cQ5f?P[=YPKTSQ7M/FfXQ@^2/^FOd#UII@V
NGXMR5S\1..54<03#J7VXY;PUB7L>JPG@8R?V>D&12D771Mcb\;K1d_B25]XN..G
WP:5)TJ:FP:@_:TDK,/X):A>&eB83QgTQ#WN642,_0CAM0[,;-4_^7N_>F5Gc]]C
@dHa#],IWZG[Q>?138::EcSL.ReRX03VQU6Xe/-Y4L<KM?YfYd_RN5L<F.I4ZLCa
C41ag8H7,=)(5;,3X]:32J[>H?.3\^@BT+H=bA#N?I?>]LF+e[[(.=64PRQgb9E/
U[CV?1;6H<=NW8([+]d6SS+b]eX=DL,HQEX>CZXZ,c+:EJT^+5&UNQY&#a8g5]dE
:_.><=#KEX9Fg^2\V]5DIOeA<FJP];>_,S(F63QAV;dFUgd8:WNJWR30N[=FAN7D
c4LR69I;H&4W4b^D&/+.e>P=CKP_.e]eQY8bL-/I98;_]H+gB:d6Z=LcL\ZE1UP1
O5b93)Mf-(H7\:PdYKF1bD1LgK26NXG>,68g(ANBNS6&#dFA8)gY42Q:@=SFDW]K
7EGe_bFSTcg0_a5gW5TY1P#E7.F5+=_YD3Jg[M#Id^ZX?&B2S#FFKfWW@ac:e615
cH#D?X\MNGUggdfX:5#Y8d;E8\F>R6I:;,(<cGf,4F\8KJYKN-N5NeA:<BB-5dGZ
Z2GJ2R)LB]Yf#@TMKM4R7g3^=X>RR5a8N__JNKGdI/baV=Da&O128G>-X_f,YG<@
?YK&74Y@N,cIYXV)-:=#a5/)?N_HI9=fTS?A75L#L)^DL;_gFB4MKJJ4_O;B)9BR
4Og/b?g?9K,;89A(?+9ALG<b?@A.#3FbHC5VGS1WGMV;6<dA60DR.;&LaXdCRC@C
<25^2d5a>)6@>e.1Q+0#&dQ3HI/+eV&,9^d,YD:Q(ZW1(@.0A0P^\X(7&T&eY&a[
8;B?3>A4H51FbPfN^7>X+DY)2fN-F-gLaQ-.=FJ4;a[<S0;(,H>RQTHVG.,:Bb:P
?(gaI\+XGT96\T#3YNEBg9&e+]2SB+NJY4(7[3g1.U\J0\-(OIQE+@K=TW/H=A50
BeBf\bNP7PHcYBL)W=KP/G\7e>?@F/:/DO)4PX([9f.3<eJO>S1aT>S/3V9I98D:
I/>\Uc<aH/B?2C.SCM,,?O]K4dM-72>W&Pf2KW6Q]\<SZM>JbK;WEWUaK9/J&.BY
R^X\594AgFabD9eR?^OT=7NYVL7,?fc4bC<W87=992R]Kb=GG<2ceZXBO/--G/IA
Q[E]00E\\2FM/),6+(^Ka>,S1?AHJTb)CRYCCL222M6f8CX8bX4U?^b(E7aWL=U/
&T3D/[?+YJ(.NNH_=.TOHe/.&CK8,E8YdE].M3U=T?_De[7LI0@I452E4_]#6P1E
)eKTYa@KT.@7BUG;5SDZJ98+Q_&/?-3^_&.T8[-<<XPI)f607)1=/WU7e)PW2I[7
&@-;DfA^IcKT#3B]_W:c]>+]daLD<Y@H4+gN&449XQ2:36bSV=J?RST++<]RA#b[
B]]dDCL8NKe-=MQFf6P,eM.dOf1//2Z;9PdB079>Z4HI/B=TZT246#OJb^1E6EVR
CbQ1AII7aLHc=XDN5f?&_H#8F/0MdZY,R_4^SaA\=),/?IMe+JWb#,GP5_d3=bC/
(E)())+;#T.,7EEc=91;8JU1>g>0QOENXUAZ.??KDg.E=@,U4^V5E7M^[bfOLeDJ
9X[F9^FZ02FgTNH55eF/LY>)6eL1WD);Y/5:JaZ^(M4EA20@H9G/T:TMUG1+I@UZ
/T_?9gR@5CDBW)O3d.Oa>33/CG#.gZ#I-eV\.gb,KDJ8G;^Vad^f:-#K=XG;Yd89
C->\I_(@eJR9H]1XHSaWCOEB)e?W&,S6HUc+3A2O]LGXYS/,YYT:F4D\X+M--JY:
9?[#?RdEP[Odd9M0\Gc=Yf8>R0GJ>OA^+/V;[0PSgPBZ+@_I;1J[WIULK#<\V(Gc
XB9]AT;WMC#W#&#EV:dN5(523-MHX25,BKVf@<^M&D:IM^dIf5bI93d+]BJQeagc
UaIXEI;V:J7&\a<b[O9=_)6Q55GM5cAC7[23P)6d:0MC\SE4fS6bG=;+#;1193\g
6(6]FfCCV\P,662fGQ(U=_>@.HOT\Je054_fU]J6>P2GJ5<9J>_#^XPJU/#cf8>[
0P2B?\@:/OX1Q;=QO/POY6bb60,&bR\U@@WLE<\Y1IWY+ZZ)Y4<053\BO^BCTdJ;
dQYVP)>(af)/;:7^d-9^5^JWP,16NUbCQ>fd>#Ea(PD(;8:^0[3d1UEATBSa^gC=
BHBF+XbS>70Jf[,L,9#\TT;0/d&-F.F<_?A[XB)_N:=YK+bPX:]5L<=XFAO]AQ:#
TfKeOQN[SIY\fTGSe63Z9,.675)5-83,M0T>NfI8=GW2b2HZ?#A&/7-AKfc;=AP+
OAbPfR>_1-Ra#&5KEOH9gHe4;KdIUBV^KX^)QW3KccRd/gadA/63K1MD9edRT,\Z
Y.S=4BS+MNVX0fa@/4W;;X7Wc8Y#>UCB-+(R9#2&g(a=EB5JQGS=O(Bf3.<Z8K]H
6\I^9.;J-RM,:Q8-+-,02HcRCR_PIFRU#9.8cM:KBHI^b7EGC+Qb:MLSGDUD360f
U3NLFDMa6;cZELd[Z5\O.)e=/=MScgK?O5LN0OTUD.CG=[d@JeB4T1H,b5J3\bE#
;c<5A4RJW@.;XVd[UFK059_W_BZTW1]P8ca2GHOI.\\D=FY>WCVWP5C_@EQ7)\&N
>/#>#He1<O6WeMc9[Cf5b\H(?e.9:g7Wa_:d?R3RaD1:,+G_6OT9YXPRfXZ(5cb:
H\5VYC0:U7[+a#S@=_Ofd,E#3cd@]5g#8g,1(XYZ?E>98INAa#P?HAP,Hf.M;95&
):UCKE5ES<-c)Og(:]W,G>H:Sc70AN-fWG&-I8b^L76WVQBa=;.9LKY]9FO-K7Z7
T@7:()[FZWe+^f,1Bg?K9R)[URACW](.YK:,O:GV9E>^SabW?9@;C+XL2(3FTgY^
@V#,ZFP/2R.X&cg1c.LQa._EC<QVBPWS+@M,?b)JeK=;@\Y@_0FYE/;Xe->C:eV#
TK,9P:NK5A?EW,ff:8,F1F,HNe1[9N09@b.>J?\<H0UNLILcQ-b3L?5B?)Ba;Q(4
C-5\E#JHLg.1d&#LBN5Hef86>a(7+fTTcQI+e6T;A]edT.+^?f4R)eg3H@RA3Da@
AXF)LIRLdK7YKXO2&RR1Vb8LIU[f2CLaU>7YXN_>c:F52Q8>X&Z299;[@6R/aI6M
4.f@?/2R^75:S^1UAC.,9XgM1@M,/Y9/)D;NE=3B)@ee-T1QSa7&,ad?>G0-^Z>2
WN8.VM/.[KT#DVE1P4/:&QPfd<@2T_T)U;f:ffaA,,N?CJ@J@\I=O=,c4D]HCdPU
6LAMSDcYD&c@Dg)0YgH&=OT/S51])@0USZDOAY6S\1G4bHUJ?O70NA8aPT44c00/
P[097/=AT0X(Z/5:+V0.6@,U.4<@CY<WAfF[RI2@/@/L#Y=CCO,-cP4Q55>>O:BA
KN76E-V.f)R19ZGe9Jefg-[c5FgIGABIH_a[9G0=K.6(M;^P3d3&TbTK+1^dO(5+
4KbQF2]DR/=9R)eg</<=b6Mb7+1,R47SMG_ETYg;6O>H/=_AUGD;,e6LJ6=d5AcB
cCQIB2?<6c;>Q.5fQQ2)U-=BVeCVU003P)M+f\bN5(CY5Fb@0J?:;1I;e?]5_,1^
(7_5Gd?-^KUAg,9cW^K,SA7Z&MG[H3g]9OgU&45=DZfeOX]b.,T_bRQbDVa<^)cL
aCGcWY7.@#]U0+6^Q;4#eKGG30M:OSb:8WE_c(+UfZDKWUN&F<S3@7#YO5gVD4])
JEOUJ8Y2b?-<#CMHfC\YcZC.Y<JZVI7CdJA=D#?M/N.W,BN#K=9D5,YgT/)#A8g(
U=^UCWT&^@bd^.>,-N.f8>YUJ1TKe-@#(;BVOb2EC&e:[FUR.bSM]E.XELLXBOgD
BS9I+W#)]#;YX&bT/b18bBX71gdSf+KL(2KHNW?T<?PFX[(;D3L]5bW_#]LXf>a6
397QU9?cBSH6-=Fb\=EcUb_Y][U](E5#@)?#1^G-GUE1=,?-EM_R]/g),DW-+#=@
=bK5=.e.:\dF8\PCHQZKT8UEXUJAUUd+7eJ.f;Sd]F=2=YI&A0/[Q0a;LAFW1S&f
)?[W(GWff]a<LPRX4?2+XPNOf&[)Lf:9AZG[JY8e0G];Q4d)K;@6,X91FPgH7WgE
0.DfVfBP#LeHKaeF@AI^G3_2HJG/J44WSUNQC9;3E8&_d0B\g1K\75^(@a(g8=-;
a_QZg\V_2+C6YQJEIFDPCJFZ\b)7/^&E:S<b4WcMB_3J26D]5XP#)5G;?M,bJ-LY
&Y-PBCa_KH6\UY55=eIb1MBP6e^e;.4c5FQ-T@K@?a5LA\,^:4a/GA,G?X_?[:CS
Hd2_TG<D/#X/<a()DYKF4?^QaBd<NQ?ABGQ1YWO]Ib6J+17Q3+[RQUE&+U49V.KZ
#f6FSIIQM#>:dOWb<:I3-7\1<LOfE6/+9;J40M.H)O/327[b^BSG,P@[_,ZD?R7/
E1Sd/Z0-]ZRgR-Qc<8S&83DJ&+e.eWfe-cg2]#ERHeAFQL;F99SZ9<ACZFKIZBX]
#]#VPIG/geC-d0\g:1ZWcabU;^DZEXW0/R3;DV-UJI=]+1&ScTN:9\J_?O)<G.R3
)HL_C9eV2M6K.cVU^?XfGc<LL_E2<Z:7(e=O^L=U-&#(Z(a(e&?7\+T,dY=<Ie_(
dTRU49Pd0\CF[[Z;6RMWC3A-bab33FLZeA7BMHFKW5La7d0dYH&]7U?/T^EBJ<#.
8TIPC&@f1;Xf>/N[>CYUX.-;)[N/U6[Q7D?Q-WLC^TBc7.AZ>J+HHdOZ4X9RV(-7
VdFB_X_FI@Y\>-[Y7\La?de(1KdHVM?ON9#H-e3\/;;IW:@JZ+cH6Z@L&)RY&94N
U_KMN]QSS3X=WNT1D2A>-AQKKgdKOg(T)d[g<X)FRLI5BQ+EB3.a4E.-ZaD/WDbU
XS^)49TFOdN&I.=Fd^+@W&G@E1E4@F.RcQ/0SH/A7CNA:XHP_-A9FF>K_[+.2#1=
-+e#8?b5.2E3_5Bgf-bOTJ;I_4_+2K(ecgY3UfCd9C+-+W8X<Y7\TWEb87Q[_B1S
I\G:C\<If;;X,G/f@,J;eK8MKGZHVP(>]Cc],QU>FFURC:L.;4/eA8fE+Ke0GKDU
N?642)AH.cIR6/(V>9,Oc/I<E4JHLeK0SJ@c@b(Oa>Ge>7;VH0KD3T@HBc>E[=P3
5QfRCV0Ee,<PbH@@S,U?JfH=YDZCJL8B_Jd#G/L+Mb)EYB);5E1\[F,26I4MFe44
4LEa^(+3(OK5NXb=GPQfJG-K&=c5@3@U#.I\K?a5U4];O;50/;QT9^M=#5#V=NfV
bJ&<&Xf(^=GN,:9FI#Y,MT<2<U[gF73F+/FPg;Z\PG3JfHUQ@\T<(@[+-agFC;Y5
Q:1b<bXH(4O,9>@ZT4IecTea=\LWRGFW@f+[+)2]A2G/F-]5bCUBCR\+EU\SJH^0
XT+NU=STa>YYQ1HA03f)g9F>G-:V^>:GR:&49[=2NF,I,U-eb],NZ8Wf?]08S5U/
EE&BIV)P@<P3L6][\?[5.P+0YJ#F:54>b=C<?=JXHN(PGcO?M\V>;90]#5LZBM/P
TI__)NXDS5d(>1^fK\,]J0DAg53/9?YB;OGS7&,A\-&_WG#)eB+)?\U/&VO)8fZ2
WW_RN87(5->X1MRJJ+1\;@?e)e>K7[5UK<VS3;c),&+3HE,1]QJ&&&fE?\YEMD]N
?L_)N)Jd^fSG7^#&MFZ._8I:1Zg234D3+)QWeF;g1U4F/7?#_gZ4&T5.TNS(\)43
MQ8:25)_YZ/FeP#;;E0LLXJ9Ld/?T;048:B+Q1dZ1F3g@_.gbRe)>,6>-d+T9BK;
TR3EOOR>^U6K<RSAPDLD?&=WI8TZa/ORXbf7D69G@DIeUJ\T+<DQ=@Z\X0LaLF,=
8gVfT^R^&gX?O0g&8-F^ea[-@5^F1OK=#]G;_2\JcgdR6)+YV^g2^,d[F,<3BBEa
FWJQ^2ADL_1CIH3N;7V40(N5^gUX-2@WKeJV5OVI]/>a,2+GYX)SgE9Ef<60(;8.
9f>c.bL0447Se@F5c[11ER1QbE5gMc1?4#g2T>Y4+B_](BZ-O\;B5F>>K=AAb=L>
6-@2#/=L@M;?EZ</\Z0)],./E6abdJ;QQ[L?,6SgcCT=^5YY+@V7d/YdbC>G-JTP
QYYKVaRb\,LIJcY48Fg1B=^K5O)5H(W/66e3-1<F(>BE(I>[S;aG^IgKD8G]?dd:
V#f1\/1bZHO,R^I#1]+1-TC?g<BN4/@W,8F@g7?6a-+&,/@PgeaB0[>6MQ46CCSg
A+JX2f?:a>[aZ3^eZ0KPDGOKAP/EQ>O+Nd_&VLW>OI#JQ.QL0\&+/)aX^LOPfWS>
[QQbFK/0,[gC1A/d[\L.<[(QM(N?O3WL39aEI:YbbHAfO\?M)5[I)G2@0KQ+YD>1
3>QD+SK1^U[-7_XQU_e)<M_I(^?T[1RUOG8TUTeOMK6RNA^=+>C=#42^O4F0C^C>
M:N_52(@O8LVOZJS-&UHcNDFO)@6PP:W:FIY(S0D0d3D2(dd^SRE?MF5M-M7@dgK
N1=-;&Z[b?F[9MUf=0\J(e9:_#e3S\?(<I>We2cVYe]<a8cZ1.C_N#deE00Tbc9?
8\X=c3g<CMUR]L>;<N?H0&_D?:fX\aX=B;#Y5[D#<Q=M6S.X3FMZdbYeNeDRI7C-
&1>.\#a22>0I]P(L.627D6P2(5IVMSO;8&OI@@>;c=LddHLOT<a]:^3)6G/]>-FX
&/-E(DM@)W^V]\D\Y;N]NQ+UQ,_81S,;34S9WS5IAXZ7ZVJVGF2:#Ya+cJ];?@Oe
:/X+]OHH+<QEF.ON//3C)Oe6(&;DHc(ac;7RN3_fY4U(_=6:PFQ:Y\KLO;Ag]8=K
)]72dMK8/:WJ-0b>R2[79=DYEe^5Q8VO#(O;5@5S53#F[6;6c[@KZC[6/T[XQMI.
bLPaFD6(G(E.R/(=Haf<-4=E7gZ4@WaeR:D1(AJ,=_eMWcO+)gY5.gD:1LeB1D0)
1,MQdgN7A[BIY[65fK-_7bF0cLaC,62f^JQ<B;a\HV0CKa3c_[BI/QLPN4g2\_W9
W\IAEQ(6@)KST;5RH1ZUG=NKK^Q_;--29]2VK(H)\UY^282K<2I?EHaQ-)c@#S>B
,S]315GS:@UJ&WIe,YJ+OI<HTIC+KF#X3563:H1,#X_,/<Ee:G1\X[=WLLR;OWRe
6M&CR[9X^[33BJgc;_PR^SDZY[0CN9.CK&X&E^97A=;HH?AIW3=aEPe2:9cH<.+A
#\fAC9B5:=bQK+H^90G4K^&/6eOQORIYf2VH[^/GF0PJU@>3UGYL-MQ0[Q,:\JT+
@OI2=2fH&V/[IM7XMY]=X<1d(TMM8)PWB?29(g5_Q9UYf-XZ9X@V+Y\E==e#?QVH
I\Z;M5,9.\[+>?0eAH(V2:8TM9NSg(LI)[XGT:eU[AK<FAJUC=fOC0[2dP+6gV=:
6Z,0eb:_fZ/>&&fEd1dbEG1.5bK79SX0H#QaF(GHB61aJf<RT#_ZfI9<GQ0CVP2?
.BBE>19Nd#@XRSUCT3:@HJ(\Fd@_,(Qf8Wf<CE.a\SRSUd/IGAP/.;W4Q]1ZLP\G
YD/NXc_C0<7[3:L/Q:HJWd4HEE;\=SZM[0SVG^bO/3KN(2=LKKT?H^8RVf1Bg][]
^3BP+7<,7VG,;IXcOV1RMDPNRU[e=fP==39+8W[RVe4^C\fB,FM9)S\R<4eX1=GS
CgUE(OM;<\NY#@S.d+#Z-Ub^,.X1@NCd=+e04QQVJA[E5KPXN==Ug_KGHD=S-8CY
,,YBP+MfV6X(Oc-HS69(BXX;CDHPWd8.^J_X#[[OPBP<V45^RK]RGJI_WG[Cb98b
(=TLJcQ]P?5fcWL-eab?4Qb0Y;2Na2G_?OLX5OF)/VERGd=FWFKE3BAOb[,1#Jee
V<JT)<[C9Cgg7P4SVU-da+G+gfJ63:R,aR>H21P[VP-D,[P]@@11?Z-WQ2F67,O0
/8)B8<,-]^Y#+I;5f+;1.J3,3R6eM8YLeC4=K<3V&UKB&2]U=<)7CHdETT\cRI8g
#fD+ag8-gCIa;N&D=-TQ[\:_2FTO,L@>53)]Jd+W,1\@-4^;2<@6\;#CHeWf2V+P
)+(P.T&&aeN\]30f2NEc#>(T@3:Q>GWL:/(G/?4R0FLU=)[ceC6+SWPQOdLV2R=<
=7X54/.,7eAeX(27&.NJ7@:7_^7&,@(CJ76/P(IMD6KB7BL<0T8/.:8d@@L:)BM2
O(aI.Z[,<#W6N_<CG+bdD?TO;UQ#+=G2\6CZQR@IH226+<dKWfRN20MC(6bQY]3Y
Wf(B8SV89IJ>^J:[G:]OdWgZ,c]CWK0L>W<)J[_EPX_;/[4&L7P1R6J4<X#3\JZf
-dQMBX6<PGAUN:,+V0,1VBJ[1cB9&1&_][c(_)UXX)TbG/[GAK;MfIH4f=V>.9Z+
N2K?M=6@T-AeIP4HA\<31GW[5K6VI<V(HM=)O,49S4#8c+[#S;X=<@aAcUCD].@a
?+./1NeW;>Y\:.0),]LF[)4f&T-d28-@\VK=54/BeNcC<gBDA22Da,.KZX/3G@\S
ARIP3.4=aM:-;(6HbJWQ-:?a3G]FN8=1g&^0E57[0K>4PZ=:KG\FH@(N4SA3HX/V
F<9N2SP>\3ON;=5H=2T1X52(<,N>?BYA\4BR8\6IHU;TB;8TA5GWJ.S8MM-^2N0;
D6G0^^2PF#EgFC4F)Y9eZ[9R_I)O;Gb[/a--#NZLJYNM2Ue@LOJQO0;=X[/1,2Kd
7QC3bd<SB6OG8@UO8YC_TQ>6@EX&(GXL>WH=La0V5;#W<J>gV?<&JeNB\8DLYLMB
GNY0gGT.&+3J(8McF10M2BHX)>Y-V5_93=JbSfZ8.[(D^.[7S4Z+KaT0B?d&-+5S
P/PgM<W:Q#eHPWROEJJ,YCCUEe^DMXBee,f#^1bUeP]>1aC7,8feX;5eDW_dZgfU
_\4Ncbf);c21/H_^YS=(c+8MP?CeFD&;(OPA@f,R&def\cd2>&T0J1T7c4,BT4<N
U<5]M2UR6R<UU6@;U\WDS0/eT4cKQ_cHF(0VFRQ5g3T&]S7E^9DTG8FU]65c(]Qd
PcJ]c5<QZEHMc&R_48,4/K_ZHEQbG=(7/ScBQ+J4;4^#.(A;aKc\,]=S:@KD5O_C
eWUQ#/M+a?XFRRM;K=ZK3@ZaZHCWRIYbPc>+2LgQbR,.;-,_OU.=-I3XfDg^<bd?
Y5V1YIJaPZS?<8UNZ[T[CHZa5$
`endprotected
endmodule