// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"
`define PATNUM 100
`define SEED 8721
`define CYCLE_TIME 9
`define DEBUG 0

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
E+ecK^[;??I9=+>3NI&<;29H:bJ:QF._?K/<fcQXGZ6bg(O,476E();OCU[P/&ea
4@c^1QO.0Y3G=RAQ91UM3XYG;eL?B\b\/#IL#5>c4XQ3R\L51FOc=fG#(ReQY;aX
W-e]<)\IQHYXLBL]C;LI/D(P&3K[ST@cWPUVZ?3gO7ef@@+/PQ=F8^EYLT047TL^
LP;G\\4gEOMLIN2&I^XX@Z+&K^d(S(+UAK3_^\_FR_.Q32XT+f2f-MH@LN+)HdFP
CK[)BN.YH[5DT&Yb3d/XLVY7X5HZ3dXYb0+/KNSI08-^g5.6:g809#UC@bLfaZ+8
J^;+8RdC7cA>3dR7LT,XEdQ3,]1Ub;IAS+LBBA_F-3QVR^NZ3E6R<cBU3WfgZ5Q_
bd3&E<V.fP9U)DHRR0U<8ef--#([[[GfUCERgG-CXVPETGEXF(Yg_HQ4F3Xc(Fc?
F[A&)6[MU-20(e_,fB2Y72YO49<\51HdGR&=)Wd.X(aKg2\ZS;K(@(+37V6WF-WG
M,:#]E,T&5HGRNEA5LU_beJ;N1N^P\YB-#?QcJ/[N]5FH,L-;A23LNUIbN#(CN6M
^4KNO\N&GRP\]F3E)3)B?.R;-^Xf,\NTG(I.QM&KgN@D.W@SB/4KQ8)cRVQG#<Wd
>^0cB\.P_42>GOIG5c5L4#dT8(g(X>QZ@C9]?@U-_53O5;)f=VRNgKJ:0(K(PIQc
WbI&F6R;O0?7AGVeJY@[Jcf03RVFGgCF@C^K3E<KKM[\[+(SR?2U;/RbDYNE/e=&
T=Y68<]0JASa]g@]2V5O.[>eA&YaeOV:P.FE+G#-9MJ<F^ZRDJcA(AfD/E^;1)Lf
T2=XUTR7=2N3+Ga/7[<;WY\bITX#46dGR2@4Zb^Ta\M+,0@.4bG2Ic80)E1JTO8T
=6(<:fY=L-:JdE)0&V,@07dNVILRLCR3aB.+aIXVW;/@gG?Y_&B/TD2bKFg+_2]=
+-7:/3f8VJ;MEgE[,eH>YDA>?.F69_USC,d6P=C]1HN0_MCL@PCTP9^H7G-11C<@
cX1?&ZM&]:aHb;0LP1Q3-dV4OW7b?JA_(\43>;)ZIc5NUWZ=J5?8/6SI_QW(4+cA
#S5T)3)87K<^P+BRC[20\NZ\c09US18gOa(RM#bI#e7ZSP7\5N;)13XeR/UL=[G+
a=dDCF(ZX:PA)fD95^TWaSQP^MLTLdCA7DW0:L7<Z(#4X1Ig5U9R4aLS&+M.65&I
R^5&)VN:[96GWUDdQ\bW5OFG1OUN_@5ND7NRF/;&ZPJQcRUU8)eGJ\:B/0&Y\fP?
9OW;KXD/N4d(P:RIdc]cI);7L67A19/I#)W5(Fc_(F=/;WM+KQMCPeQE4)DLd4cU
HT3][@7c?#O;.S;-;4e62LS=E66b3U-eC=fF-.B3V[LD\OP4[_::?YB#Q3ZQeE4T
OR>M3I+HNEL=,:657J.2151[7Tf.e=BXOc3&BbaN?fCJa-)&HWXHe@b@JEBN@P.a
g<QdKe5^#QY;dZgDX4Y5KT=7C#.VN@(5eU8?g;Qa0N8Y:>cU?+9\TIKf=R:<&cOS
UW+5OKUQ]+U+I/\HEfd2@cB5H_L#]f&3)S05#?-9D:UUFCO\M:7WCHR4(7N9L;Wb
R_262Xf;87-8dMc/bcV:4/@K?QM.^d5d\,C:fe2,dY#B_M&GZ<;,7X?_\&OKPL6X
(=F030.-BEcHXY-gg<0P-UWIPa);QN.FgU<+gc8g&@;TRX?e0VIS0:CWK0[C&Jf&
+7BR8)\4Q-5@KZ<=OcB@\Ce3\TZP(E,;J>73:G,Jc&bGW+FZBP[N6@R^A;5@KUY6
Va05BYg_4).<;\,bE\&<I@#?^DUZK_)U;_>2<Td9N-A(S5Q)YZ=PF6d;W@[K@Rdc
)VI<FOZLX_?6,S?-)b4#3\ZASE<0O9cUQBV9)<F(1_ALeeL2?.-LfJVN7P7&T=)7
Vf5UKL,B^=dB0[\NSU[bLXJ6(6e]fELEJ#cM2M007_E3ecB+.Q3?A<Q[#(Z0I;>B
fc+](Y43Y[B1O]/b@&71>Y_0<d-<I1Mb3)7VO3?_GF>J_JaNUC-C?M;.WP9#F7TS
HNbcS<@9X/>21<#3T9Q70,MRN9<K/VSSda_&(bN(3&YZ>-3.f6L:aKPWb5d8[_-0
R=a_/&dJ:TQHS(dH_e].;Q=cSZ\bI(/,^6UI&O<e,]-H97?9H1][Tf4a@^[>Q-P,
VWCbP?1NX):R8EfER+B5RSNRb-[-QN3^@6<4<<4^db8>5UL5\&OHGc+0I>Q9B6Y7
_9YK,Af.X.:6UB-:=@;ZgNg/1J<f3d=BO&+6MK]eS>O+-?+Qg+GY5IgQ)&D<K]T0
Y^H@HJ85e)Bd^BXY1AGCN6MJYR@fIRTAbO5Ve@gGdF8:e.@:EW5V-@.TAf_cNBa<
WG<KVL@@/,<8P\X/E71VgG/8FK1XH(?(eHFKW/Q^OE]5@.<(beTQ)[?[B&3(ODT(
ON26;W4/COXgcR)@0<@R)<M@Y[WK,@Y@aXQ=@^^3K-(NZUIA>e<gGd4[@3@?@Z68
4^J+TZOASI6FHgLfP<NPG?N,),1JO_FRIV/>IM0OI=bg\G8(XS:WCdIe+CSCVRXT
7\:#AWUI#8e.8_UK+F7bX<BS[N_3B;bH<576gFf=7V[c]#f5F<:&U\I=TRbD;X\E
g8SG?@,I9-0#F[GO<^]DUeaAO6B91FABYD^5W2MQ,-8e\]FT-BGe,;=0_Q@<XWc;
33C.GM)0E1fJGOA;7V@RZE1d2]L(QP/<Ff@_PDNLV;FS6CaCc@H=96FB@H=F1ag2
9SaePP4^G(0ddV7D:JYQ+eeL1[,gJA1NOT+TZ.cQBHKB#6<0^[NUSTf1QPSDPU4N
F^_Q<c5C3QW1]O@.&g[>4c60;&9D?88F]T_O:<RXL>06@X=b3=eJX^/4TG_(e,(,
.c)I#_-CKIN)TSLVI<WR0=T=@B:[Z6\KP3OeCYH3W3T/(a<e@ffT___B=IZVZ9=@
O?6.<+Y8aF=.(G.aSK5baGQ[8JNEAP6R4AJA.8d6LX?DZag9.1c^</R7B_^\g,e7
W,@/V?P4OS=3aV))M4+[MQHXbD@0<^aGEG^U8Y/7U35E^[DXGb<E)YcLSL\d[_^b
]FP_eHQB,a,ESV)@g/<0=O,IB]XU77Z>c:b@FX9ZAO52:c\d4Me#;J[_/M7=EY&N
6<TX_9F4TYWOJ;TV_V_WA^7TS8[TcNS2P-GW9bZGMG:UHSXN01?_S]T,;6<@)/M<
bW]-&d,P&:VZW]b&gXcV4)a@[:d8Vd/D584fbPO9,H=@V_(64<b)Q@N/[=1H&4cL
8=^R6G#82Uf=[)@U9U1.D8#<(R][D=C>OAU>>\4U4<OPR#2VO=HGK)C=.3?S.MgN
UNAcVDXgWeM=e#^HJUD-g:;:Z?BQ^caXFg+9(AeZgP09;M.g>6ZQa1U<TNJ7_aXe
<E7I6[N[[;6Ggb^Zdc\aVA/-\L5T_78-c9RVJ.5G9),(+\6SI/M.H=5HgYX-=NE:
1?Q1^>T^-M7KZ4G^F._76E5Q0R0\P:ZgJO5H=e,B941FE6E/6.]P8c7925B3S?47
Jf17<7b^L3OA[K1UUQN,H7LQ14(H./@S#UT?BYM.8QbURb->YD17Qdd+eH_99QD<
OP9NU0[?62>7G_QHVE_Y9C]XFKcCaFLJ.]1K4NM4I^BXP;UH_Nf;.HQ9[,/,PU;V
J&HL]=e6@O7)D\B,+88+c]6FQ0ee@(S]g_ZO.F=)Hf3\XH?BG]AK,EF:E+Ge+.Nc
8c1N[Bca8.a40HdAH^7/adLGUXJ#(G;<:@TFC&\4O(d#Z2?<ODNMQ:7.?/WZ=eE#
f^L95g^X\ELWUa-WYC&8_;=-a;>YQSD(5+A>e]&R0eUC67YeD+0V3)O=Se#@dM-7
Ja:<GFLB+Tb@9)V^FgYQLC0#HTNHO77aZ#-J^H4)DT?T&0,0d?X/U6IU64:P]FfJ
>-)DZ7cE5[597g:b/G[\Lf:4CCN]GQPDU\fR(X:I)e,?V[F\ZEG\1d2,&N2bP8>=
K61GP+^G>=,]\.I+aTWG\=?G8:<YOV3?/Xe1_:H6YbC+\35H:)>SNNF[8>7XN2RJ
:6MVCGC1N]bfO,=##5RUUUedCJ5E)8Ed9L:WBf1R<+^V]D9^LL8\\-TT[fYHe#Mc
ZDSNTG\+4E[,=Wb.aG0I[AQSEOd>>(WSXcZ\P8,ZVBQ==R2K<,Z,739^T:OgC:ET
4_:Z\]4JOY^N?WCGP]PC,2Vc]b&KZ8[,P^Od(>=&VJZ=AaZe?Y3(XSNVVV\XE/3J
&T)WIDOKMB)e6P43.^5:f-#^XQ)F.7?DPM:XNB+2c(R&0G3BNc?YSaXK]e@E=?a6
S&2JARFC?M0@(g((@BdD2]@#\E(#:#3.\RZ_dIR0P^:\T5NBf^&2a/S#XHc7ZNP0
YH&3<]]==Z^<L0cOc2ZV-dWBPJTOS6:?4;MZdaL3g88D_[Wa_7Y_+0O_8M]&)bH&
K\-]Da/&HXB[]=+.CgPM?9/OES;_3_Y+2A.Y04#,&_3aI:8OHH/P5&cT,,f))@5A
@1LH;3Q=DX_I7,^3?0bO^X7UH;LT(@I+W7R/=+^6eWF#;FUU6AC@f>KGD1INYE;=
:GHAV#S:KHB1R8TbY&.CII3<S?EMBaUXb5TfZO,-:N3EV[@GBM3D9[8,2&aKe4@+
FMCaWG;(HbJUZF]JVUc+]Z:ZL008:B6I]eb]aZ@.GQ)=ADYM&FMLUW3g&Z7#_E,4
9R:;gRCA1g,WX2>B-CYXN_4(XLg3a/9F^?d48],YI-#&g#_[L8P(7fAB]H)39P3G
KP+EE06Fb83646-5@302]S2LI^UIUQZ),XYF@[KM\KRG;=?Z)JO&(d1KdEB>FZ87
4U:FG=>#YL5fTP#PJ:VC1[gQM=?eVQ0XXEG#cDXLL>\VM[2SDYY7Z.<MJ=Z?VM)[
TQYcEg/L\X#@?f5d\,^.1gXD#CEcM4FAcPYcO=,R(@d-#.:?<dXcdeIKe?RbPe?e
M9696<(\/E^b&3dc[bGZXY(e)[C@L,3(c=E-C;b<I:GWfO.WX04N&/H0JSTEdSD&
NHd.Vca/7>JL^4.b)f\fN#6,E.CQ+DX6?#7]6-CR<\6?Q\KZG2)8-)-OLQYd>)Bf
a#VeJF/b>,Cc+@cZ?:.2^VN8XROGG4fFGeRY7A,.R0#4.gX=BCX8;e0P>gHRdg^T
0=IH=eJQX+=J)WQMH/KONTAU-caY9W@FcH^_7M2:].IL,G--3P<W]<A5GGgZ3gb:
^e(GD1eKN;[RK^bMb\LP12=IJ53&[/=8@\_FM[,[C;L_:XLa?fBb..aWU3b?CCdQ
TA##b0\Dg+7cWB072]WRKP,1FU[=@bD./:DTc/UQ.7-TLTaIKE^c8=W,OY:1O-a;
^,c^cZ&X=N_aV#;_g2NEeH9O9#.6QR]:3BIJa<^_?#Y4f02,N9@.&ON]c,4X1;1S
UG\<W[2cIEI07-Z,0A5cB5>D\[8@<fKD.7S<SUA2(2f1NIXUX<GK+3>MGIT/MAKd
-bK^:eQ,cKOQ0f6H^TL.AgTR?5@>QG9/RS<6BQ6W[gOBNDZcKZ\eU2PObN4gA8OF
YUMCNVXBLb^Vb5-GGIJ?I117+6fWGRb0MTW2#WN^Bc9?30A0Ac-O^9CS&SS+^EV@
#F(2aBT(gVC-)#=_<P&b5=J2#,QX[-;)<F09I<3\/YV6+=K<U96@A\[-d\0P=\(e
QI>2A.Z2G_?9#-)ebF0KZ##&0bS\UX#aX1IZ5K_@f4dK&V=JJ=eQ#<HZRU[\eOQ8
[2#BdgS;^QKFHa96ZKQ,d9AGGa-TO7^DUA-C-gK]EW]a?eOM^a3fU(?[/A+a]gGV
I@A6GOF)Y3PNU?A4IZ.BNVH[//E89+_/?BGHJd-T+>b<=ba5DM@GbSMe+bWNXf93
P,aIBFB3bIC.9Ce4NAB91VJSf5>Ff_MM(TT[5H]1T6YFNS3>YaXAV,S@5/U@[1W^
YG9<^YG)Bfd)I[Y^;C?C,?+5.&EC[2N5:Z9=0gYaeHdUG.L-@L;NK/ZQ<S),dUgM
[NF3M_UUD51e[a5P3)/]c?5<A5VU&A\_cQB];KXC<0?_X8+eV3ZRE/F.;dD+gS(&
9=eOFP[=O9T\K1=]\N>P2AI:,ILaWe+\2c\:6Z;CM^JTUQU]MJ>dYLVf4?Q,G.9I
V-bOD3+#B8T@aN?X.g1(7/TB\[R^EO7)ES@g?)BT\#GZ==IgU7J=>:Rc([PTC-A(
-]YCT8+6Ue0cTYI3gL[TW\WJ[H;43WDQT+2/KBB<]cI<X7a(OXE157(^S:/).AK4
FW1b?J5BN<>P6:MXG-)BEU1I(1FL\&:XRYJV2X5V3(@97^ecODaNc&KVWTY.KY?c
RFH9E\J+O-eL<\AVU&(EEN@b>PFd\Z\IRE&T4]4b?:,3)fP)@XFW9eZ_3cP8-@a=
];KQTL,e)A/BIfH8M1(QQX(>S7<Y6;U@B0_@/_e]K7EPc(TQ.LJL2O7D5W?X4^[<
OR,(R>,&/G<:3IE;5&6aB@A>^X5d;@N5g=bN;W\F:X0EbM:@Y?Nee_+4AD<,RT3I
K]8]+<XUAO,,^@JHKV_Q]-C_IOZSOT,2@[^HPE50,)&0HE9Bf[I>RVF?D1[CcP:B
94eM/0JK&D@;0>J?0d2HV7O3f]&4g&M=1U=1.6(IA2Dg3KTa4Z-dPa?GFQS5:6G\
YeBY?Lf)N>ES]a.ABL,J)5C)X88M[0NC=KV[QH>=:#B/I.M#+?:#5,,U?C/0bO<@
eI<5+ZVd[Ne.E)gN3T<FFM<c;2cVTE^M(H3>MQIRCbPG@D8/DR<1U1g\WQNF:f^V
,S0WW5J^OM6a5SD:8[&6_HWd;TGR+5D.#6c1^bN]9/+3Q)Kd1NRAcHf3>O1>eZdO
bE\-d;eQ_C52VBKYITb1WZf&+W>:RaMO]>1VdZeJaO_5P3PYO<;+YWFT?_/(]e77
H,45S]]\#eJX;:g)BDAJe7U+DQX_W7f[F;#)Q7aVGRVWK/KcSa3.5PJB9#),7>Aa
\KX/KMH29[^?K_SFXC6NTgKQd(bM4KHZGNQ5/=6BQ\^Nd;3.9FG]2JUGVSENMKfK
1._IW+=ILO6[EJK^0M9g7=/RAf>>-<J8-HE0.c1,eSKUI;Z)N5L\ML#F]M]6a@?N
)Ge</^:FB]7Z.1>_U92[+)]:?\\KGJB_c3?/OaN[S9Gc</7#K_H[e_X(-ZLROQ[-
SMR+CSd([+N>dSS#^@-^6LY1EJYQ=:OgB),<=)&/cHQKJ+G8LKAP-TZ:D(d3d9R&
5,cZRT+^P+S5#5-.8_d:D\da3<(4M..,5_R5KC,1e;EEQE1-E<7Q73ZCSUUdO<22
U-N:H3XJdc\/OI>RA@W@E)#fL<H).ASdDV)2\)Z:T\;@>1VDPa=N_:522RNYBZO3
7QM_eGU3ABY^YGe&K+c@A3RcdC_a.HI/#1K1(f.UK]VOOR6GOgO#F8VK5(;aW95X
2e6M[_#)>0?)]02e=4T=)A_\BdNDZB&,)SbI8(Y\T]-JBNJ#gT7NT?18d;V<N>ZJ
9EOB3QNgGJMJF6,@73?FA@M;f-ZGaU4Z0(N)@4IO==H\Y1+3#_eU],@/T8;M)cOR
RMB@TE6eIg,B\D5-Pg2E1YLM-<;XLI]dMW7^L-GV-=?0\2?,KPP:P51WO5_3.AI?
,dNQNYfK7;-QMW&^_MP@d(K63GM<Ha5d/5Bd1g-?;4b2[)O/EUS9Ia<[eFNJJbRH
0.aA3U.M1<Wd+NDJF=eR[ZVeV#\+Pfa?2c^I+/1c0NUS]FLBY6V8WHHe:G\.+gB^
#\E931Y;Vf^VR22F=2OMBLAX)?^ARIWOg,\^cPE,gW.3Ve;76=[+4/3;;8+1bGJO
JAW&1ZB\_bN<\:3bJMf^b/9(NS8S<[1adPS[_2F-&Z@_ARdB(P_OV\f7=RcW2V_V
KOI#O&?SWQQ(]SeI\US(E9+PO.^E/d.&>#cLe#.\(RX:XVE3QWP;R:Jdg\7f-Ud)
F1.VSb.EcDNe:B17)K[=1W?8JCDCD^a49+-1=34+g#]SW=8D(WIKad\b=KaIdYfG
0,T3#=./M_ZM,KQY(@8a<S>@PF0>&FcZ1?g()eFVJ]:1KcGdOc^gRE+J&<cZ,R=a
3AB>XK;9eCZ6TR3e3[5Cc28MM,3g1/?(M]+aIN^M91O7X](b62(@)WEF_\.7g[&I
X<Q1eI?gd;SH<QD3>)@[eOT:f1#8:K_29fIegZa6E5I<(Ie.P2-SMD7W^^GBSN(6
3ER#TI;>38&L?A(IR,)e23Hg-)59>HYJ2=6K6F>]L-X9T;F5ZR9QfAS;NN8ZL6GR
(N)60Wa:0XL4M8ZM;Pa_WMTE]fB8RYf#2_W>9g8Xfa+D9Pe1;<_c+H)fL)K+Q>A6
8dg9e;(3CMX=Q<CF(+5M4SJH9^Z[NZT+\256C3daD25\Bf^OGXH7agW4dYZL0G)5
Z)U00?@fbFeCDNW[GN<8d_IKQW/AL#JL9B_5bYB.8G;6F<E7?I0H)YTVNM/JK_Ub
C-+PNKc[CIVHO6Maa,#7/?=.^aY[e9D(9P,e?YW(cTbAPJdgeUaR/R_(;;P,O0f/
QG/Ha(^^,BLU9^9=N5DP4CbHQH)b<bJVBP(9b6TK9WXAF0I?4_dQ;3D9N_N1LAR3
aR-JaZZ#HWg.Ob:86b(9aE9If<G-,aI>=8ZMEPfVfVc;A#I[TV5,AWV\-]E2e&;Q
KNSW<+T&+GAVY;.^:7XIB4[D#<[\Zc7Y.;O,N2ARO\1Od;EUM&HF)J?FT7N?M2I+
GLf:/:c38b#S,@2JUD>Y5^DP3])<;c5-+YM/4Ac5Xd,@?396;P&EMW6MWALSb7CE
Q;2T7bcCMYdQZ>/>5CRQCGB5;/@Fba(?#.@EB?HVT=-fV^^7cRWI<Hb+@E,Q0C7M
#ERBV9_M&2aBf;U/X(0\L4f;)L+LL3dX=HGU(U1ANZU6Ka]5I+<OL:O,eM:<@g7)
(U[M83;^W&:N\)7)]P?c6.NfB,F]R,@N)=SB).98B24L,632OP=d/;AgS<2(XL(^
\Q:HG5@cb60?RH0c9]=EbdKD)+Zd:)>TYcHS<=36M+N=#U1P2N9>(7UF7OY]c,8H
dI>>0#gI9^e6O=fg:;E-fD-7;;cB6U_O)R>19ODOOJ,L.Y#832&b;,_fS?R0UR7]
BPA^WQ\a?YT9(fTPJ/2JePHP<CP80[,3fd>:+.]G(9EG9)dWDg\GPF@YSR+US.YX
IJ<<L<>Bc7^LMX]Z,-7R3D:F^L:EVSI:<P74Z\<Q&@JG2fdB0MbOb\S[7#BGA(HI
C@VMP1GA@TO<PVBgIE^I3)5LAJ_0DVK(D#(H39#_TO-&??RBQfd2B:.DU-#NdOT;
I)RG6#bM3SMF[K4E5]N,d#DBF+(^SaV#7((cg?;<8ZTAb/Kff?Z=RKBWMA8W,MRB
X<D7FQ-\^MecJ1XP-TNZg0K[2c(@&0.RHM765HWMB5=5<4[PO^TOZ:#MU)OUN&/Q
4\a:^f9U\HDM1fDAMSTQAH:a13@b7B-=NFP(I-8dOgC&PINT,SN9AHAS/TI^cY2]
Ne@fObIe/S;D=3J7@[XJAO1_NbR.PW<Eee#3:FGBI7X+XCQdFNbJQYS&3]fOgC5)
]cF2A39Ub@^^dG#Ube,^MIL/G8SXAP=W1W<JP/P7Z7V7;W,2U\S9)Xg#]&W4N2@a
247Y3DZ6N<G.6#)2V@5:AVa,.&>Jc(M[cR;B]?^&dL8a3F\+G7FCX8A#_BFKJU@=
<Q]I[[(^D[fKUZ<EWJbU&+_1aG<5>8:DD9T.cefJBE9GNe;f#d1I[&5^@\[+Ub+M
^LG&A1^bC_bF75f8:CBX;#IY2d]JbGSdYUc9N#&9d:<.RQ@V;3]FP5,+QLL[HcE<
Afe^GP1gcc<OXGG)c\eM0AW&E(<LK.A0eW0f2W\3eY47XY:;\FYc(U9[-K]9CNN;
:bBK]_G\S5HB1:I;<e/a[8GQID5H5U/<:B:<_^B4=gKZ;>>#G)U73T370O.UOSM2
O2BK(@5e:BE;/&CZO&O39IQQXRO.JXG<^SE<NZFgSGQaU(F(:?E+9(7Z?JHF90)G
C_&2(_JT;W0YI_HC8VK,\OMF^,U^IY.Y3LF>R+V38HWGZT3>HHO>dIG]38>ANgfE
B,9L7^fLgCT^8@N?S>PL/8@cOUcWNBf:[)GPB1IVZGV7-2DF1]5V(OSNKT(8-=ZU
D,,KEQd(ZV(5b4D&:U/[T,eeQ+#ECHK:+MYGNS8NV6JF&+XR)CQW#;I02QX(&L]H
?7B_#A-)NT-F9QLZ/.L0KI/PW2-I&LdT3,&5#3;433ZdCeJ&M9fI;MT0?<78b]<H
PK:WN_=^5+bKKf]^G9N^cY-@?KU#B=8CK]Y1=eJcQNb65.Gf_&]^3_)NH1O<:SGY
=PDNOT.+eE7@<P9a);G?@+D]DfBBCBA[c/6<U4L#XL<D+.gNN^+:+fNC24eI2(FK
f^3>9PX?CFLO5^78^1;G:b2X>)A-cY:Sb550SSD#K16MbQf@bZ2cJ>]O:J[Z=<9V
DCe>3TPYUW&7\WP1VEdVJ(-FTONO@9eKB=:8L1c+CI8aPMc@\gJT?N&+3c_GN\Xg
TL7a96:9Z5@L:O3HSZX/#2&[J0HS_O3+I1U&3)S8K1Of4Jg]&aUUg01]d+[0P77+
.,U<[eg8-@Z1,>]e0KG(^NT?;KEU0b0KeUc,J9.Oa0)6Cg+D3e_FV8(0JbAQ:7C,
#5f(aNTcc1+UHID=0<:f6A>V/TSbO.9KaY4F\#U_dEE,;CE.8Qa^aH^PE7:D4.ZM
&a+3O(KI>Re.6=Ygc&=E]8f^5]\d[\4X0bXL6[\/=RB/GIH)97&IT@>:(].=#bc2
1=/+2J(T__LD:ZaEUKJI80>F-^,RXO^^VC]DU3]XV@Z^I0<&R<=fTaS3&RRVRdE]
(XO.b_=<g2^HN?VW1#PS>O4&McPZ2Z<fQN);JHL75>GS&OE>8DIM7f_H6b8Z[E<>
14XON.5POH[C92TZM9eOcafS5[TFP(34M2,2Da-M&Sc)CBNf&?Jg4N[?[0FNR.Ig
c1;4Z+B[fAe(#]ET/]5LD=+JbCN:8,TT&+6F\Qb-QUOU[M6<GB++WcSD&/c1Hd)F
)(F9f?(.ZWT1T1HJ(5P)bR/:LXYEA9F=<VB/bDKe1S[TNTM@K\Y6,&RZgIRSDCXU
U&<4]_[A_3&43]&/_e>A<Be@+LIQLd.g)2b8KLLP-K\R-NfLDXa0L,&0OEDA,P)D
PaPSR-1:9<1?Cd99JIE_VI-Gc-S./2W:PVb6^YKdcXb:dcGV,U0&Q],[=fV^@^<8
SL5&cZD2f:eaK5Yd2+eAaG?.ZR[AHS4Z4,dPF;0Pg?gQa^9MA>386^aMISQD;W8A
BBFC.\&7(#b8c\]Zf<6O4&A)b2:VNFO[DI#^/FQ?\?A8JSC4E1M6O\0_]]9EQR+g
I^<Ad:5<2^R9^5ZfJNKSYDMX0T\+f+;^0I]e(V:Cg?Sc<CY0G#)D/#S):^adO>?_
c7dSJI)#:R9.:#.3G42;VJ,C:SB8c0F5-V<g;?+P\4>]7a97PF#6Q)Df=QDcc8<+
O&U4>A(-7&8d,[P\CR#g8Z[95G@(,1]^C=7=1>E2L&&)KD_50@:8PcD3:B4a>WU]
.AD5=bOf\[V[OI0X,Ff>RAaAY&^6F#Z3(-\<);b(8I&b#0RJa5-8XI[OUR+5A/^R
NL+/DV;\G-1Wf@133-T(FXWE4R+4&./PEIRPf>XCJ[-J7(9FQNJ3NLSSJ]@M.>&1
5fNH&@\B+96NJS\3YS?2A&Y,/a9>?98)>^I??F;)MWSSOfDQHJ\P@d[3+6OG-e@B
Zd,1K_Y7_I7,HbMLbV^F?:7W(1OcCLE>)78T&P;cYcUE&f]K&4JREMdWA0I9V2VX
>[c<aY/,YP\S^AF4#gXg79c37UUH4.XX:_)SY[A[WKCD(R)afXKW>FPL1+a#CZ.W
F(De@_a\,D8dZ8c@P(2egD]\#;4d.T^-R49R5I<b081>;X<#dgHW4Z2<LAKC101b
EPJNLAGKQS#\#ce-RXY+W?P/X>bF_50Q0>]GP@BIH[a?4&OV4.)9YbD&CWUeKcI:
3VOYaXI6^^2N@?4+ZNfG8F,95@4TYJ<=3)G?5,::N\X0&.F+T4DRO(4.MHM02_P+
QW>\YMTF&:QPOV\&ZU3IK2NW0PRF;FOCTG]C,NOcgF<QY7:\bcd9#S4&fXbD_P;E
J#LK6K@N=36S/7/B4a;b6;;ScXC>a00>N^aLPbgUO6?NgT#Xc9;UHX8;NSF)BFV6
O-+@b#RV/VdD]6YYCIT.INEaD>PK7LQ=a?[<Q\\,AP&^IVY4W7]N6OPa3^&7.QBf
C=MR4[SKQG+gM(-UbRZbSU72/J?2=MW+W#ObdAQ7&NXR1I7A+LDeB3([C_\)+&05
5:fO9I/;#>d6/442LFO41QHZS_HgWK<9RQ0BE&^L)TAEBN5.;f-49d0#F+9gQ.dD
Wg]-RXW(4W_VD)?4LTDS\)#<:9cB@b<,gUVE[X[0]J7D>?5V4IcaO-GdY?fIT(=Q
6V0Z]A=VW(fL#C6d394XYIbPe<40XMU;<OS(-V@4X<VS0,f^g58:Z9(U4,)([+J9
]L8);)C:,7d6W?5OO?)C4\dZ^FN5N[UEABK8GSSRS];:K_b,D(XE4/B[MR(Q974V
A0(_42e031aUCOZeZZUB/)K:aNB=2JZ68YX\HZ=QOV]Vg9+cJ[[][cE)WWYbD)a_
]/_7Y.TV</,4bCN&Ve:914TEVO=L)]Va1<;FGHVd^6Za:[JR-/(5S3E,N[FA)>O]
.cB](AHB-e]/_ag)Q@eTGSSF#&W=#<g=L2=?Fc?A35/QG(G0WEV)D@^>NU]^aQ8=
/]J6@9,0L.GSQ[J@(_R(3KM,&gF1>XTMCO4:V3F-\X:^NIHVga[13/H?EHXAQ^/8
:F.DKJ8W\58ITB1ZbN(OVf>&RF<PJ,IE/Z)8P75RRgX1cJF05:,&dVT2N:E(3dQE
RZ3Y0[dVWQ?+;7/Td2#Y9Z657QG0?\M/;UD=@Z<T5@=]<V.AFBX\gCH-)G<?N<b<
&^,fB<6TTOd?/9;LE/7gJ4WgW1O=CJYX/d9ZbU+g=91951ZJ@=^TM-O6d[a(LG/P
aL1SUW@XJ<>f7(A)1[RMQ>6FTTIWA7KREQ1PGK7LSQf4FFNX>T\QI-+?a-DFJaM>
F8_MT2+ZaJ08)+bB[-NVT3>PVg,JG3MF7(0:&[H_DQEae&NI_)KfRf)ZeS#P]EH\
P:36JG;<;<7U?:R^3@1gK@Jd74[U55g7T]@9W/N@,QZg]8;(B12WD,(FI)c_61<W
M@[:Yg3YX)Va\.KeJ3/[/-Pd-BC=)6K@OC&);GV=de=]DQ)EOQ.gg/EP^XE)Z[\\
&GQFZ?G3VFT4<(7,cL2QUNeJ;D1J@2;Z?;AOOA;9)0aF:=,E>?/d&F4)a,g/HX-Z
=6]/dcARe^8b1I=<B3+2E3(JN[Q)da(USM[>8JB1@/c(f:3WZ[9.O2FY.O;e9f\\
<HNa^Q_/9XG+)T?IGGXTC:UP9\)>4)0-UQ@^;:_fOcQIbXEVJ+Y1[-MGN.?;&:B6
HPK0#,CbgbK66PE4W5>A5bWb_/K-:YKEcO)UAUAA1F.LQJAQ=-51@K7,L_GL=fHe
P2D&FAWG5=6,.GD1/I\0K@.WC],-K7:Je20c>Z\/Y&O/+_S5@IY&,KO1=L\H+GVS
ZU+LE?Z/bPb[E3gONXO7:MR\fZUAe7#MAG-XBKb;DFQ^dY#5\L:SP00US.L5^3Tf
<He5:,>>W&#c^QEIZL:#f6dXa]H_P>S7dB=,KQC/TRT>2U^A#88b?_>.(BKE#<5K
-M4B0RC.Q>VgK(X]X00#Of?=Q7N@/N>T\#X[^X]VXK>d\#]/=^EAW^DSK>B(D<Q-
J]]f-K/D3SgDSFG91AB2.D3ATH0L)D=LNVTd3;U@98BZ<<3IUE?Z41HM^8#9fOJ9
]HOT>_E[e#D&-gO9,ceH9MQA2UA,LQ4W704-dSC=aY;BSg5(2U::=1_C#3=)EYA8
1[@f^=4AUTRT:WVYgFHg?#?4Y=T.Hc2C(@:GQA7TX(L^8G+KNAP2_N^6]]c>VYHL
Ddb^^#FOfGE1VeQ;GLd:IL(Z?a:g^g0RS<RK)cPXLSJD[[F4d[Z4VO+dJB7#+29M
DJ_UJWSc\9CV[fNOc6N[05Qa3@5C[U@7/>:c??6Gc/X-)84X,YT.D[5QY:HX9&<[
<0&WUFT]ZU-\9OSf#g7\;5/C?\M^R++[OU>TV0<Ag+]EI/\b9DGHQK5M\E<YX],8
^>-&aCSQ#M)CYc8d8\AacP-&-9>SRfW@Q5\1LPI0H;(1N7_V>-[(,0.KVRfW84]c
_RKN-9f>?UUL=P=(/(C96=dU#X@PDd)Ff@J<aFD+_+8X4PaM&\Jf-O2Z<>0,OD5-
)PPT>8\S11LRf\b:054.(0\_>]^R@A5-:SD+^H@S:XNO-YTG4ZR@gbcU,Q^BeF.1
33\ET+W+,-Q//94G>C0^J)H<WEgXfdRcI/YP/V(N8Ua3K,C3[=b8/e#c1a=H[>KI
;I,R3BJ-,]JG7DBg/B@3EJ2D+&U3Fc(=bTb)<F:?_7PL=]F+b<>T;0F=CX&03H@V
L5TMO</AHE77cSTFZUQXb5>,aHg^X(cCZ&IN2Q=IY_#2b0FY-6C=I0,S97,fL<fM
>EE1;MHW^^DLYaa^.3db6c,Lb,[CE6(aETAJN/N08,;LPfWYH=_d^AE^Uc-D.G5c
acA5<XeJe=\/#^P\a^2_B(\Yg_8\5JdX@cKU+K@PRC8QcED8@-9TB\#C._+e\X,H
8RQ^5WSSJBQ41Acb_R#DFIUbC\RA8dDSQO0AJ+#X33Mb\KJedK_W?+O(EPP/T;.9
C1Q)G9W1NFN9N)GO]HTQV_-C/QK/QdMUV,f,0YG+;8)BbeDYW_ZYZOZJEM^+L<S5
.H0?&Q^\+T.0;7>^XM(IFNBZ@PL.[=)ZUEGDd07ZeEb#OR[0&f]bb<:O&HL;YJ_c
T[EeA#T&XQd0#e8AR=Sd1bBQ,b6gc726I]5c@</E]]@&V()L0-4=KEQHTaF&M3&2
0f59BC@0c85T7DDX2(YaSTF9cHX7,0]#I)D)a-JBcWcF1WR.7aT:(Y@@(4-P[M3E
Z]KT1BO.P1KM,ZGZbXM@;@_OSG=,V)WI4.JY/F:2V-#,dHa=]g.<XHLHV8\0NbL;
f5_UJV(<5II[SC^/K\[gPEbc;PP0@_I?NMDe;?1Y76BPC)dIB.)cG<3<_5)cXRVM
N+T0K?.a(O2?,LgWRY4CaS&K(ML7.DYB@(f6^V6OS,T^X(KYW7>)PBGV7b9A6>,f
S#e[^J<2Q99/O6AR&:d79\-+Ba;G^=.6/+[L=JWN7d0^_\fFCWdB4]Wd+?PAS@Gd
A&Z+MP_I?/G9I\?g2aGKC2G.b:.T<bbNY?@e[<(8L9=F,2@U&a,@U)B5Y/K9:YHG
G4+e8SJg8a-#MO99+g7GS:SG3>@)TaB)[@O&^(&[>5/\:+C(+HMZG.&#I/L6@IaG
B8Sg+SeV&:4d5:@K]8RM;#47+7[J[f-96J/Q#O_5FbB0HWcOg=+a(.N7W/+TGS^e
4&@dg?./QT(ZGUD<E9<\+2NPNb7ZEVPC)275QU5_5Q,gNdD5N]c7)Gef2>I2)6^<
/CQc1ZW>f):BOTWd=RUL7L)P7g.EcG/Ka<d_W&JLA\F2f2SWa-6XbU/TU-GbG/]d
VL_ANS2JMbND0-V,/EIN)V<M\P^@?OZH\ZXM/EdHOZ/9\(J15@D-=))A@9fCI55U
@45+b?^c_0R@01e:[T>2f^\;Q2Bb^dJCVBBH1ZVgXPREfH^6b6NaA3Q?WO?Z=^/;
UL2=^9bHUQ^3@-P2g-HFC1d]cWGeY_?)]RF8G8>,d?e9NALF+P(&)eXCfaZ@d<3A
f92,BLB6)SCY[Y?@FU^\1/]SF4R>&E;0AF\7Y<eTRQXHRYXV/&6#<ZeDL^SDg<A:
E;;Oa#,RTI#MLD1Z9)BEd08dRP9,DX;9Ic6Be&7Tb-Hg9AQ7fbc6dUL#BRK=e-FG
bcGS]<[IGc=dSLR><X@H:<O\cPMIMWL11YMA>)/0<HBC<Y\#<JfI+Q+/4^<OOF1C
B3XV#10A,-6WY.aRf3P;,ILRG&AfO>CRPV0eKc[b+e8e61@eF_U=9W[7c00&./dd
/<3b4JCJOQ4#3)3FS0)P[/Z1AaL.L;/IMKE]#;#P[;Y9WeG?S(VfM&7HOf6E4SUC
5.XN4[fK\d^.8F[)?/R70d5:dTWA)X>^KK64UcR?I^5O08H(5-H08BdgaG?.H.JY
.5gV[dTNUT2=ZXdDf.3aaU=g1V\PK7fG.5E^aI:\7?.e[_:>XGVPH@HN>YLDJc6@
/HT\UU7Y&cUUJ[]@Z7Tb]KX09MAL0]IOS,6NN7IA@b)\2#R3Oc3\ZH-C:2<f?WZ7
TK6S08M85+HH.:HU(g<EL#Oe@M1,Q.,\/EZ:2H9F-g_c>H>A37aeb8E&\+dGT01e
N5fDf)N\ZTY&f3-]+Y)B,I6Y(&d?@ALAU8)X-0;KFJRE(#I@]EX,#)(-;dXXRAXT
S3B6RNUTW+1_J(1ZFDXP:\AF16UVNJ1)6Y-F^g.e#b4P6-]NUJR@)VA5[]5U<<gX
<,?@/BO1eCgB59Q?cEU<g,[e<GG;b_]?42AWHf.=cQ^J(L@1&7[06-J+RQ;7:Y_V
7L8OKI0fg[YFc1W>PTXK5b/STd4FX=>KH11HK,\L&V9\C/90XK]):b:a(dCF\<K<
^g=7[9M-CFe>Ba>^D=^_K78I\P:U0LKC3d6g5Taf^=^RMMH4JKV(I(PF8^N7Wa5C
c6FTN7LXWD5,OdUgE-c9Lf#E<Z=G#L?JeLgN0N_A?\>JIca580WV7.YXJ3e21HC.
2<1.>HbO9V^-G^cC:[YD&CTMR]N^,N][,1<8Q(1=AXX.72D5/cVW8N6/(QD[W>Hb
aJ0+/72g/[L.VC&Ra:Ua]YE6Cg@f7gDa,(+@?/44SP[8SCKgU4K;1eI)-,R,e_Y8
4G0(E)c^CT]DXB,,NC7EcV_H[,3GST9)>+e8+EdA5,X39?FG@A07#2[.UWd:+:Lb
6R;;dO3L\9X.aX1bF.QV#_-4:PQWW#Me^;O<b2S.ZENXcTEN0DeZC;cL(]&K__)]
/Oba)bXgCSLT95+OI;)@b_@WE\Y\5We\XL/Xa=&@fV]_)Q?02@K@GUfVgTY+bSSc
[K.<+Q:,;^Z:5KJATcQCWA9C-7CSOWVQL=f3DY]Y7Q_XX9E=d3&RVE@5UZIN-FfX
6d-N_QB6Q?VC/:=VPGPG,Bbf<O^&1_K-]ID_GAR^-/8F#a8@+,bZPNe&)CKe=C7C
BCXdBW[EAC2FX8CBC+.A@4+,^X8^@1]:2CQ\Ra?V5fQ;:9Qf9GKFG#a;=L288ZU4
#[5,6G-c1@N?6MXMEd[8]/JbYN.OYfX<AC)QPd8HJ/G^?4[a9fK1?eda.>d9_,Y-
.#d;IUaDEAR>Q2<)@&#_,BZF2E[BTT&X;Q\I4#=@-Kd5^JKf,+)O6T9R1>^HGL,K
g[X#)OfT&gC)Z\8W1bV,S?7_Y/8^\6E_LWIDN,e:NC5_01ROb1NSK/\=D<fdWbH_
b?-daAY_L=MY&3X?/&H2a5C,6e,:fWT\G+(d;fI6NZEI1g\TJYU93>&72V4O=be4
Q<\W<bM@_&FKX;(O,dGK(Q+VfW-OI@T9-eTO+NZ=Q_O7&CR]&@IfXQRg#&,.-TZ1
DH6Z)bO]e=M6Q[]-:WOLf\@T>,AY7^ScMdY8?,].3WOW@K;C+[:D&dMBe:&T?+[^
2&/2VcXE<@dfb3,Kg@<3\Ug];g1@4g8E.c=gUA\Td5W:a2=17JCY\-BU^S)/&(C]
=,QM.5WT?=K6]C9Y6@#\7BR_4ND:YDG<=Pe7??+-]UY=BM@F;M8_Y#[,aD6?>K8;
=b62(Rdc/W-b[P+TI@W.P/?2-PdDgc=DfS\Q>C20]B:\51J(Y@6aaKfHZ.f1W;H&
E:/-R[;)PU9B9;L_g2]IF>)MX8V#W?;/AX^DHS1)&C0U(BbX2@/+(@=.[C2:;NPP
Q]+J=RK)PdT7Q;7\TVGDB39FL?Y@g#S<@Q/aDfc1[\E-H2SL-9DGggHEUC,8[49M
91aGIC+S(Y2[SIX>+.T&X;E7.RZFO33@;2PV=A&)XOO/_g91JPQg1LdeFEC9bFZ7
8&K-=TZgC3aP)-(.:,4:2CeDB)Q0N>#,UF^CB0#-M?)3.M9#a0>KP;W;@JX?3(33
0U>fL0+gZd1\GP)_dK&W038ccU895)GNZI#I3@QDGc]6VWN8-MN3/81?Y[CafMW?
b8+S7NL:2UHKKY_c@EA^R=^:fD3Ae3#_1-B9MeW0gYe+1(b\/O\F&M(WDB[_Aa9Z
HgL\7[+4Z;L;#H4OJgUW))]c(A9O.&C(^AZ(8R(E(>.JT;beDE?FW&T0dKWKNe/0
T@4T+De45C.RC?=e>.GD<F=_^Sf5VWQFNMN1B^\4&7]:^^D^I079d#eK47@62#4:
Db](Nd+3V4K&N.gN@MVQegL5;<MUD@C/]J4/>I3^-1T,PG4/G];<<RXVBM8<dOZ;
.aZfLSAB+_2K0[JVVWJbg-/b[?DeI.^UJAgZG+3[5SFM8P\)82/X6LT4B/H@6^dB
Seg0,H?;@&KLYf&LQ<QFC4OGSM8@5bW&@S<NS2b_Bb1L/f^,BR&LH&B&f>cL80>3
X6#g+?/_ER\Y(=?0(K1=.@4YSJ+L.0#c)M>B9:OG76S?23E#Re=;=GC+6\<+]U@-
JLG#B]CK#U3c]XC/-4ZCDCbfL=3f_]/\^?0fB4a&DJFAaX0X]dg>b2/NaO:fNB8\
6H^(,:e@6+Q/RDe,Ve,g88@_-O.@JL)/BYPA4;9/S:G2KF=K1ORd:?MO#O;EWg6I
?Zf-32:#6LG9WfXLD17,D;<HbB\\K_S]6(M=bMbD>bBDY58U:XUbMBf6dVRE/6>K
^.O&^0O5495#4?_2<U<(U:CRa?d+dAae+PL._d0#0e624P24.\_;XBe2c@g&)X\;
:@9@3N(]#-UFZD7(>VUNSHVg@c8SN\>E[_A&c<a(9D9HGF7QM?I1;d+g?dPR;a8a
.AR>FgB?/Y[Z)TUL>,Wb+GKISN3KNg,Hf7]5Tf4>M5d&O@dH/EETA@R8LZ]2ICXH
7I52#5]_=AO#fUedL)E@C1BHa11^\U(XC,:GgCWZ6T1G)DDYfX-cNgRR3Lc:VK]2
gI;aJ^T:4_MeGb;cZ-aeG+)_e]D-WSAc&.0g+X2I;E&H546_O;MU@J5DV9FA^:MQ
&E6=-JSRNb,_a>TAN[ZZDR<OGcaBOP)V[S,LZI>TA1CCR?4g\dVFIYCYX9V3W2a>
0MOOb]<=5bBD[[5ZA^0U#A\_F+=;VSV<P&)=7Cc[1L#I?I5?(&d3&V\3?&_&IeYC
,XAW1Z=H3KF\^(O>?;0YF,:^b5E3b&O)[X,#0YT/;([4cS]C&;NUQ?)^TH#_>Q45
(WT@Y(?/)g3?^1=Oda.1f@^L(V6>@5.gSbBg]9c^KJ;I1LMQ);dNEWb^&G-eM;>I
-R?f+[Z@H0bb0,759edKX1BE8Eb@Mg(dSM./3RD,)NE:bA1/S:WF@O[a_Q@M@PV6
@fK4g9X<1Ra5(/@GFHCD=8#]LT@=g,&b]\?,0+IJbP_;-X_2F3P/;U.,+f\Nd->#
[ddZfMcOPONMY+V0@,T/JPE#Y<Y>\dgd5f/K@0=gTL_3V8[V^+YfbJH&K<C/Q)/A
J<(^[/)F7e\IX\aY:VK0aGT-,2QJVV;SSV&RP:2X^Z.5^^1HR^fM2^0Z=f(.1=O<
g(R>gPMA>UCdKJ<D]b>0RcMP1N0_:74:#e7Vf7/bS?BU:A)[B[D=P&/NO0@L.+&b
0KHJ[F#CDZ[DT7X8_ML;?MG)4+&G:\Oa#3T;&MERN>SS]DJ4GGQ)EHeJKT(E2O54
Laf8\5G5AY[OK+X#e,T:A1PfKVa?.)FV3O7OJL-cReJ(W-aaIKB+X/LKC@6&5.)/
-0Z7#1[cgG4QPdeaN<0>W_R>58Ed:)5F(ECIOP06?Jc.>c>gBK556G7Rb\6B#&CQ
g:NF?X]F3X+)>eY_QE\A(?Y^NdE<>246GS?7]C4#BEGZaWKD-#6N&CN_I]-+K@=(
,S7X<-/ZE48#D40_\g=1e]O2UF<-5D=H7F^)U];3TOa1VP3.B;>JF3MA2AdH&W</
GS#)c\)EYL&/Q1-g/+P1CKHAHX9]-c3NR7D5/P^NM#RI[_3[aY=aEH_[ENGeM&<:
\O,bc,F7-H.BKTZR[([)#7JG1^VR8_XS&;LYZN/]>.A8WRa1=SN,Q>VA1H1/<.MJ
85d]06dL.eMG8F2S61dM6^cgU\ZV7?cJ<MKfV<3KYa_+)8aM4JE-+_#&Ge@Q7/K]
K]>7:YN&HV>,HO[;T?U:?KK?Z.g[_\ROXTEU_SK?a7(KPSSZcg+HUZRNXP.=2<,S
VK,JG8&IH)cKUE?,YL+J1@&3#W_.e97ab7SH[bN/Vd&F2?3(eWaNJ9D[(O;GCCR\
:.[HMYF=Ufg]E>#J37\PF9^#GU+:8:d)AZ3J>6e;SUUMC@?ZbC(461H@QUANRE)U
)5@)0QP]27E6UKG+Q3S(HYIQ&)>3=gCcb.QaXI_c@BRW@RD::?N8,_;+))S4c_K)
3?A<.=g9P.?@J?M[U#baU[8O>LZW86?_?E:<<Wc]:4a)Q4EM?EgeEQOFQS35H<::
Q&D8#YP4JK>:&^,a7[ON&_0g?2-Q;YD\R98&=f]:C\,L6GSCZWe3SO[3GKS#-[V>
cWW;U:_E,4b?16(H.8MX4P(FHM\0L&:9\+.7bWJES9]PIMZHUSK6N0]OeLIUYRJ_
_0R9#^CASXON0(d14S65\e?[EH\AV+-B>.RUIB,:0Ld+:/#0D=6/IX@?03AM4M9+
SQA6#8RQ4U10=&S_B&<gBb2]O>QV,\\0:Q-Y6VR,@ON5PZ>Cf0>7g8]7.SFH,b(.
>[D(+/9)Q()fR98XYVR:/OT+AJG-=RW>HYg7H#M6#d(M/(RFG;&S#;X=&XOF>T8-
]=gG3UGE)C=dBS^@N).E,997c+(X5b#72d_&3R/FK6&FQa[V,KQ7gE_2];\bB,Ag
7R2VB=TbI>2V=]BaSZf0I)A9dZFd-AS3a7FN3W]?3fG7Z#<QdQ,Y=#J3e\S-,R0c
;^(/JVO(&1+\80.L(ceR3M/6eIA]X4;41_a#=cV.MJ693+D#2DB-_C>M9S[d>EcG
+O>UL-c\)@g/SEGBJJa6X^>=50Ha=R[\IAQeg-aHZCZ=6_VK<F0?&2,V8_@NI5e?
@eb[1\\Fd4cSLU@D^GFT9<_6+5f0a7LD-Y6?8I:EfJ?T/Q-_)A=IPAMeLTFE\;CG
5S])d-8P._(8_M(TF)HaX/71J#=fd=T@4Y&R^W33?&YaS?LXebFR3/d[=,8OeEWU
FMabK#aYRZYb69FR6dB>)1:@M+dg.I.NO3@N>d2XAcK?&8Q6&CU2)ZMdZS5C2U7G
V8c9OA9^L@+aJc-J.:N.gQQPb6,:3;_:E)N\;R<U^(f7S/RCNPL,B@-VLgaI8+_a
R30&@f9D377X59IRDO(M)fPF8D<+M;<+O/6MIbAQ@_Pc0(_)\GX8/3MT]?;ZVaAX
8J#5>Z:YQ.Dc,NQ47JdfZ&;>NV;2<JY4ZH6\,C^_19TRM1FcD4[HU+ZCMg>_L_-e
0ScI;[5Y0a71Xd9ge32Q9:EO.3f302[aU-73T>DM4]?Jc.C_cU-dQA(^S8[GZ0S1
+[eWP;-LXS>V5TbV1@BH#/(V:8b-8?6>YS]PZ<g8fLR4^85+&G0OU3f1MaI\\-8?
-,V@(7G])g<N?-C5N>;252VbT[3B^R(bO=FD[a##73OMRe8-3/9<5ZU4#fC)+WZ0
[,<SI4^PM;]WGOX)@1gVLD<0QXR(?],[/)>L33AgZ3^4AL?fT=]9/W;&GXB2fMQT
W0RKV#]-+WI[G?Fd,I_S(1<G82(_3e071;YFCGa,4b4Sb;KP)\Z[G.VG1764[BgN
;1VgNWa>T2OU]VMY(?(>RbF^(D^\O6:T,>U4A/(,3QcTP_N5F/gdK28??#Q+F1P?
AE+#PV&Q@#MZaMgL<fPHI.aK@+JJ,Ob>9\:2=RDg><dG]-3Y\MFfK>LHO&G3V8XC
-c5/3K0,O^N7Se4M?Cg_H3/J:PX[NV,[5OeY^QNI0dHOfLJ&V351_7Q,L.J@Xc&K
C0@bR-b^ROB)a-1J>7eB4Q(.\4SQSB51F:_&(d/f_gS:&B:cS<N[MKf^<@NUA.R0
?<]bOEG2&d5ag;\MAW;6PXRQB=g#O1-[]AIN<8UF8\B9D+Yf)Y+WSHDMTRN#eS.(
UTL4F?/:BB);R\2fa,O=0IU(M@2dcF#aBaV9J,bU6W##V8X0LS4:2#bd=@D-[)RL
REHJ5.,(@_RcK(d>b</)B8(Z8<B7G^R4dCIe^(G1RE;7B+V]99^,N#P_K8M8)_K=
6,b2-D^.#0X+T?\3b.(U2Qg)T?O2aeG>.,+=6CF#V@CMH++T3e>Q=fe\=5A5L6W;
J=A<[,D-OP[]5;.+(TE6+#(JCP7;,YdGPBcCCPIDG]&^I>)/#0b?TJ?V,A]g<9RF
^ZCR3VgA_a+]Y6SBfFbM&UOZZ=MBg>c7F?c5X+W&^O,VIa8>_<8R/Od_+U37)@ge
PZ80SaG;@68463[C(33B]cJ\\P=G\9SUaS04d-:=.B23)U41Ve\CP[gedHK-^(56
OIMDRR+UdUFZ@4=H2NBSWUd4Y/J)5e#Za>]#_^&_D\SAeNWa.[ZTFT+K^1L&W5S.
@=dGNB00e2EQY5>_d@a#-+>4D373:dR+MIeKU6DF>G?>GSe(Eb,_BOE-4G5GQH^A
]-QMU)=WCJ&^\055b(DW01).LQKQCN:M.8Z4R@[?Z[UMJ2EAA1Z\O6JbS1GW/^F5
e,ZS1:S25f/Ed#=AEg:F7B:2SH=@U14CdB)I68Z+?LfG2?K0WPEYNg0.EbH9]6<2
aAFSAKJT@U/<MS:QX3NRO^5XJ(<&_7+M2\4+Gff^U])9R@F+d1/\KJRe4b3X54<f
gW+=.Mg8(OC;)858YWa:O?#3c>?bQ3>8ZT/DLBff[)^/a.Ub=Xd-4N3D:##XUbf:
.@6Z,aJUT]>Q;L9;R:UDV=/O(3;M/P:DL\YN#7>T:15]KRYCK\^>UG13=15^)TT<
>8UJbDa;TK<:HEJ#SMK1IA76,:I#2,9;.;0&YBR3?\6GWc0^EP5P6e3ae,#_BGYN
BP;?dATRSL6BJWMf/C/6<,9#51CALRS\fPZ4<KS0H8BZ+d\S?T2+=&J_F\+1XDE@
\<]gMR/K5Bb=R?-04.bUVR0Q@PbK@Za<R=Jb)QA[[a:57]B27g;B954QDADQCEZG
aA\<.]#7>>>L?33c]f-\gUeK?]G#_S\4,L[c_gL:63\]gT4_VMT;BX1+F;Kb3:ee
1+6LHg:LBd]76;8]g,?&&;3Hec>f??e7[96I3><4I4\=V@J[N\X.P3b<1V]&8/0f
<e5A26KcQMe)7Y_f8+GQ:@gJ/8#>IDgKWN\(eT#IaU?I6U<DcGDe),]BW(/AM<3_
XKI)d)WN0Z.He0:^.47SUD#Zb2X3\[NKcgS-..HAf;(XD?3I]a10g;)QfTE1L(EA
/:f(BZ1gP;#Qa_@VXf[J-abCDU+[>#:]&+.QeVG5?N5CLdc.#[=CW1K)dW4(#&&+
g04.??3b<=9LR,D.c4C<)E:<\=+(()R3BE<A^7d]BTD:9.&2a7<A(>f+#QU2X(Hd
G7Z<g(>PV]W;b9&.CDGaHbg-J(&RfRA,+VK6_,GfIF-=AIHLDL-7X=b27:aKMC35
#NaN4=JE_3W6,<LMP7QKFZ+;U+6JV1+N;gbMKV9]UTJeTF#WD+8^ATT)[ENRS)?M
I<&@SYE;[.>=J?3OT9PWIgPUfN7cW<gYLa-;\9Je1++X=#=7JNTgW?)J:7eM@VIP
/4(AAE&7ZM[8UKS@,9.,9:5&BH&Q4d1C08??>3G@N&F@gTM-XEeO59/5.#8C;H/J
?Y967#H2P2-E3\_L0fbP(U(B&\cO,)^KO.S6DX2g:X-00L_3AEa[c[-TZD<+]C^J
=e<I>B(BBTb=Q_HDCP6CHPJK=b[T;U+</#B#4Q8Q#<0O);Y5=.LNXP(/cN7)62#K
>b6)RGRW93A??Ga[f2\^g+,[2C0=^>f;-bR0N5KO&aF4,Q(J&RZcf:LFR2TUE(/(
@>B2gK&0_Gb00Ac2g4fN;c=b5PY#7RI<VWM^_fMY81XL32F2(1QL.E=@bNJ4&e_^
XMH/[-Vg2^7U\,B,\)OX/G+RW<]9PAD;1_5,/>S1#,gOc/(]&YA&)3&aDP/0]^.>
A82=59QEM=\<]_g?J/)c3YSV+@fgYBEc\\2f#;2<aBD&W@C6CI,YeENT4L?O:Q,@
#VBWc-0/S(#V872Q=47aNO@H,?32&<+8Pc\41+cTUNWER?K)6IR&Q/S-KTSB6RJd
T,O_4??WSRg9S#EfLd\:FP1WXAX@@2#;PKU\TP\6YEQH7_WMO1P#g,NJV;WY<KR_
g,@,bf=Pd&DR+I[F/:&615[^#d3E,\Kb#aO:</G[PU?0RYd2\CC@IXTb6W1cL29#
6,/Z_W;6_IPIML508ZNcd?OTQ6UGg5??O9IB_?EQgFV]-=(QGIJDBgBK4,WW-5gb
WO<bO0/]]+.>e:]6_c#9DISSIR&dY<OZ5fX3-]Vd-?ZO1a]6)d&<4^?+[+1dB]#_
Y(N,BMeQLc7fJ?d]>]G&@+.AEB-I+L_DKTf17eeU?6F,5DH.2(NATdDVeFCCcbe4
&>FBTXE74G\\dZ<U<\TC0].DY1U/(F.WMH\ICG->IceD3MaKLCBN,@IT:cD=NOWf
S^)HD_JD[bc(JWB/2MZXAX\G?0-3X8I+-gD?f_G8P]Z-WBE8_L\]Nc.-6?;\0(?9
Y3Va7]P-T[[VL/)?G;,V5A8OJ3KSE[U<bGE#]IN/8g96F9U4a(CN9\H@>0fP@CaX
52c?II2RFbN:3:&:KFR)WQG]EEMCO_Na;N=CJ>-X2/J#O&;6PU:+f\aME2CR2BSR
QDV4VF#^b2J2?KSfOCB&F9AbWQOEG#:#&aF_&NR;Le2=P26A&ge/_G4[a1a(X663
Afd(TJX;G\B(P]@SH[a9IM=ZBCY-^-67ZT>8Fd_FZ&edASgX],e)O6@N]@P3P0@Y
bWN=K6-KXA4.)9D-9PH(CGg6We?].M_7P&>V&W8+<V)VP?Hc/&D/)HTH9IV/DZST
PG3#3XS7Tee[>g/J9fR&<U4GY?eM3+^ab)0d_]#/N_70W05?E<FZ]CYd>15A];];
7R?&9MYO8T37:.-B3dfJSKPS8;\NW>1/F/:.H0FKDcD;0+,T&)&(3JgE_0G-NV86
U2g<fcR^L;7D6VT:81/KT=#b[U:2;B/8gJ6GbFJ&5LT9A^c=+=I2LX[0KCD+I3,g
^]HU.b):2P^D5E/27LF2UO02?,M9(-E6<N?K/\/P&V/8PEM^0R_^4.bK^.,8Uac7
>NTYQBL#CR4LEfD422Jg=R84Y@g(I_6>8O&bU^[@FPW>5(g\MDN_CG],Pc38KVCX
+VQfYdL-1;6U98_X#;@J8\Xfc8>.T;U7?05J8-BL:R->++_Af=c@4dfQ1eVX6P6=
e=Z5Ua<-P/Sc\WQCRbQGc2A+TS?]1R00]cfXS3ZX3B-LU\?P=Gb)7T32-R6@A</7
g2gd+HOE>_57SSA]\6NPBabN:>IRG82,CTcY3CRLTY6QO2,[O:<>,A5(cV[J&FNV
).KEdWEXf>-C8Xb:dP?&eeL)TE0C@TRS>A2N<-&^\OB+PZ<]F:([)V&4B,EcDfM,
#,dbLFR1Hde>:]2.EE_N^JDR+<?;2=^0e[4cG:)J4cX].g=2&7A++fK8O9KA9EG+
/_12PHNEY#[>Ff\EL2=KL\IF=\<gGQ^F.V8>HLT.7UeN@#WFaTC[Y>A40g[MV.HG
[;]2H>\.6]T]N6>A[KA8;QO0(<C1J=^=QR[V-_SX?)L_MZg6dD99QfS/#9::?_GS
>6FaU@Q\0Z@AZ17K]V692df?##dP+@1G+G;Ug#LJ54LeU(6VBC&+O0EZ5YZ:LVGN
g6(8W@\QEbYH[,29RDfM^gL5K,Re#S\[M.a^?Y0?47b7gFN?)V&fY^O@CV@2H](g
CaL-]_BXb+CEIG@R+-JI5IER)a75Oe.[AS-2D@/.A;GH-H(#6P/RV+0HN3J>a7I4
Y1R@]FRR.;aR\]@H>C-W9Jg596dA.,[#OU+N7(K[A\;UMR^#>O>3=/XD,=-Y2a=P
#Sfc63\b5F-;#)I9@NA;Q=/USV;9[_\B_c091&A_0P>HOCXZ1IdZK6GH(4.GNf7#
f&J&61LK;OOR<9U?e.A^=PY.S_C0JGO46E&@GFCG-_W/-_/9\MHX;PXVHC[.E.\1
=M#8V9;;DF511#3e/C+VTV0fJbS??VXE:a)OEHQR=2U56a+92EK[R:ZTW1]Y9\:W
.0g:SU>b]\+&E641NEH+dZg[.(Ge_c,)KY?4eAe[0VIYZWWE3#,[Pa3TP&EU3Z.5
C:>D&CQV4[Jd;X@HcH0cL54Z.RAG0^.f#+KY\,0)TEM&fY,H<e6K]6B/1JQQ,TKU
Pgg>PRD<8dQ@f#S5=U7-6CH0AG/C2R\\]&D<\5GPR@HH&9J=JUS/dG8LWb(-RF[G
/RRNHgKY]-+I2>g#T9LW78XZ02I6(SBQ5UK0c6,9+LA&Ef7dJSP5:UQ48&.K8e?;
O)5e1T#9DUg0BHQe\3]C4_S)DU=Jg.]M1ON:>b_<L7#Q&G>ZJ;K=#ZV\@/F2-79R
T&bSaCX0C^CL1?fS9=F<GOW^F0E5-I?320^KE^WJ9WJ\]U(a-Y;=?K&=<+O0gT]P
>5]EA_>N905f?Z?LFK+RXfL:b<S/S2P@bO#OQEI:8N:/aAUe#84SJD);QXCE-7L-
/O?4M=^:JU)1OTORZ<78:6Re4A>1bMQ>Wcc/GZ)2Lc(=SSV#A>,=fNIFeBK>D;7.
N1gO;RA#=@5BTPgKV=ZbE=c:>\JV_F)2A-Mg\LPV^c69[3BdS9V8D<.:4RgT8f\b
PXAUYZ<_gb;SA66/Se&VOB<5HF251()U]J^=RgN+(EEY55g.-H/,D99L5R\ZCMN3
Vc?]:Lg2)[O2@ebb\+9:,,ZLF@WV.<YJQS4&053?c2MXddW;?\f:1d_+MWR,aZ([
\B__S/DU_bY[bcL?NLJ<&0MPI,OTK64K>\5#]1c:9d/;f^V>AJ+[W-f;TD/C[N0^
])XCJZ(2F]>MLbX-F=CWX^MFZ4X7L^fVVSI5WAV-H)0,:+R1JbW\@90+[24<YCb;
3S8Z0V#ZbJ,S:/CbR#P#[JPC)[#V<4#NDN/,--#+\f5de]=c7+,T\Y(5BIMLEgEZ
ab+.1_GfH=N.-B^F(Hf>=XO(:f+a2O@:,e+fM-3P,_Ic_L\S=HT>;+bE:1bD[T#G
Vce/-5BI4O@_OfCYV8F1Y-R_WdNK3LS/^O76OO[S>f/UBA,bX_:&EF,V&WV)N&R]
df)fRHRY4E)a/@=7\f/2W6TW@\<2<[P6W21bVH[&=+Y?3d\^dWQ=?AF#)_8C7OfH
34fX^f/DAS)7=/.g)[8=54e/b#S7cf,X,O6S\5I5V4L+b0_bPI9FRB9/F#[VYd+f
H6PgW,)/O7eXBDX_M1-0M&>?)FG]4(@@Ia./OLO;2R4LW.RIAP:4dP@GBd2:.?<@
3KXT/;OPe&QQJTWUP(-;]3feD[@_(=^>=VO2\Q?[QH9(CR4?BT^MbL9@=B^#SN\@
DM<5VXH#ICcF>f5O,)YXMEZP^=eZ?I=475IHRWLB0?OI^Y>b?G_:#G0YUT69MXR8
7>Y;JD\@_XFME>D\(>@:)<_&>5]B@I0S-[,^I1RNTaI.[FNX4D,F]FJE9-:f>AQ(
,fO7U\V>+K:C<[L=1.b\a8)#@/Jg,/4TGZ.A+6NAe-TbARED[W?9Y5/Kc4:g:EAX
<QRVSK\.W4H1R?_ZTF<@22XL-^X(NR\>;\ED&^AV\UR^O91FJLePA#ZSCLRa,#d1
))#IaKPD3QE:&5NWf_8UICX?R.?.?-8S\HI)fIOXP-Y8/>T1>SW>A)LbC\ZW?IOL
ZN?Z/0\S8,F:WW:&8B.4NH;e.4ZI(.Nb#dMZGPgca1d;7_D95?W;2N,P-b6\]#K/
(N_6JL/fIFP@1a79<9&8b>L:U9d(MD&E1SP./X31P5EDfKA/):_8.6d.WMA<2>NF
gL:6/@=>E2:6JR.(#d_IdZ+2&3)QSbS#bJg,GMa[DGX\04Z\S+V5A>).V?b-7g57
)00I1[32Yd?WJKXeLKIY9;7(U@S>J^b=;:Rf.UeIbRIQZB]<cKS)QgbIQ?68,P56
YZ>G;FP4[4A9X=\IPK2LX)RdU=<ZVNDOF]R=Q-@^+AJdM8:&B>_b0#KTVZGP^5//
Z8W)1=N5S@CU,bbTGZeC-g0(J=G=;O9B)DQWN)H;SQRI_42U/1)N,a#K&C9\U-B=
EELZ;0A30Jc&AcT&ZX^X;D5SCLQ,&L@LN(,Z_N1D)7@J7P0X_1UaLUI-K(MPQHHJ
P?f.03AR^C)+3FQg-(_#^POY-4RIM[Re0V:=G_WdAB2&g:&F=S:cXK?GZ@C>90=7
<R@LZIFaHH9ZSIZ=0Y,F+W#J+N^JU=gZ2ec,O+-gZ5>.\.H<>9NN9Qg+[^2M?UJJ
95;Q(7S063UG:8WfQ270VG=g#<1.+HN6^fY[Ub<+EOV7PAF+1?c01d/,V9)^7cZC
MT[U20KAZ5?UJ[WJ,@DBR8KGD_5D6-\D2#0L6+Ib<5[CJSU;;D:FD6A1RP.O]4D0
Z[:d9eHD4K/<ATd+H;caS#M?Z@dIR)bd8]aDM:J>Q+TTPB47#Z#-4G>0&EB#W)T>
T5CJedD6K(QH7d98eE1C3:<;f]S924IL[L0(DA;>FSHT9.4NS(;#KTJ7&Q?<AW:9
Q_/E>79T?:59+\2XJZPSNb#P6>94#[.U\O+B+.A728g=Lb]4M3DdII7E@]XQ(FcQ
/UYHKc5B[C0&^+Mc,B)9H4-B_FE:6E\B]A\]QG\8.aKBObLWV/.LBJO@_F.;>RF/
=AQOg^DE]ZD6:+0;]#4e+J1eMBHf=R4_Z:D\]D1HJNC9>f?[b.gb=Y3/ZbD]_<N)
Q8dd92+_?3+2HZWJ?\V+MKVHG@N6#LI\4fTb5D;YR/P^R^fUKQ^d],I310&L?EU/
?:B@:2c@9\F64a-,8a<#P>H\?[.XAUERA3#\PfKa<H^,7+=H2[a126M(8CI_BM_0
0^1N4\9=B3dDf3B4VD<eUBL())QHBW1\?AcAP1/Z.bWUf-IaNf0LMR6<1#]SU3N,
N^ecbdLDd6=3@c5QK&]]Q-I0.<4D?dZI0R]+0(,f9b2B>E_YD4R;^M66,]E4P8@\
-bG/E_=3)AAAd_g)PYgJ7TPKMKD3Te6NJg+A@?6&K\RJNcO3C&7dBO)==?\M@L@:
#D9&8=_#a8>X78CPg1N/)PUgR-1g47bgX(Q2_bIX<O8aOTNJD=I<f;b;\EOU@G-c
0[AMP>9/MC=C->bR9+d]0\Gc/=NPg1O;e>=NPbXc=?2T5DA8ceRePB5]3,-K84g9
FKR?I6Z,VY0R,76&7HbWB=UHKYX7BFC^/@K#;IG^B(7O(VcUUPa;M-ZM+6R[==Hc
9RL=5c35.aaB[dX4SRX_cKHAKg+O[dLSF^7J.]HIbR/0PPP8cF)9<7I0AR@+c=4<
B9dCWX533)W>OQObYE;eEeU,/LQ#K=0dN\fF0L9_+++c;\:RSXEW7gVcB^3SSTcD
755NcYbGX]NZJNg4)d7</EF4K;P,[J_7G@<-\aI8=;;MP/?J/g_C;)#PQ@GLb^8f
/g.X86bT+OJUIS_=W\f<3GRFICJE+F,HTTaH50N]?1aDXcN5S6JeME_L6B,/IdIN
S9[Ng?VNI4<87U?Ha68B<F5OI,geF-bD[<-RD)W9JMC<U#;^@ff_2EW/<geAa#eS
&,ZFe.AQ:#AO)>YR_^R=dSQLbC8032Q(QCKBVG03@KX28C/\5GCMC.1Z1aJ)/dR\
#53@P/REB9b=a=_Ic[]5K0[/g_GL8>X#+WY-,Ff>(#UgaOe=(+P-\\&J8ITX@B^:
dcc^HRgSa&;?YQgI(L7\1D]-]EM@dHL2J7bKSb(eY8.<ScUYOfe7V:WQ6^P8SE\+
O#A4A9TF)dBAFZ+&:LX?CCNU7T6N[^fKS^,R-P_7D-E@FLDOJX8&eI5XWP@V+?KS
c0I6PIU5H>R8^W3G&TIH4a9b_NZL(fD+=+]UU5I,IHG[8-/;-Sd<TdCUcCOg^TD?
JS?,1C/IW;=G+4a1(QR2cF&AY,INg]J#<DcNM.YI>>V?FS;EHI?feK#]B.X/;C=;
]^#DW@AYZ]TVL,=3>P-&6f3+6YCFKD\K5L;]1Ga5TL#L2-D>#I(_[T5H_K#X<_1K
#3Z.4TENGNQ5^1ecS.E;O_8W^d&Zd^9+8,A>:A\)LgPJ+S?=c.Cd[MDgIBRJ],A2
KJ@_^]TfYWW93NMa5T_L+Yg-4;2#f\EZ]/:ZbAB2S2d=aB7(ad3BGBHdKUc?8>JT
5#Q=-g175c@?:dVVb27XD[)M2EBZJT/(9KMEf\)8P8RZ_7,9M^+N58D2BSNR84._
af\^.-O&CIT,5&C[E\Ea3ge#//+dWIeE_&C+39V3E,f/2e8MdUGMU<)-EXZ@^97f
8feF66^d?[38B<,\D9HD=25TLL71?V8cEGLZgTDQ/Q\U7R5IYJN_20:PWFEa<f3I
D/fa;aJXA1-g5[:LdTMDXE922g7?#fL?b^6+6+&@;XU#ONI-fR@/Sg05(1=5+QP;
M_#b8=-,]&b#4UUcCC0257@VBBSbQ4#4HJH+FN):BVeX_A0RCD\U)2HPG,.TWK,/
9J+3?d/[f-@03;cc][7.FG>F\;8Z6AVU54U/d#WYKH-(/JAe@dV=e8E0/1fc[b=R
&TMP2^OWd/g;_[/)C\>LI)6a@C7>A/6d9&9@5.\R-XAW1LCcGEK\cL0Jda4Q47c=
SD/#Q,\@d^^aAVF;U1Oge2I[BTDK;+d#+cB,RGGE4/Z?gI53D,11\fX[:(R^^@(+
gIaEc6KKe>/=0Oef1-^?91[RGc]T-;+@1#R5<O15XE=6&>[aM:a8W675E^\<YfVN
^LEaZ(2H;3,B/_4X?RKc]PW[2#Ied3>BIbXf^]TM<KD+837PE:0HM9W[aEJc01Eg
.>TI&;Q1E_;RB/>b1dbKbHZRb[bU;<\Ad[@K57O1;H/H0A-UAWg,I5c.8Eg+?JI@
8:KC7&2gB4#+E#JQ^L3BM=<Uf:-2FWG_I:(c4HN_7eM_5N>TNYd2TNI8@R?a^0T0
WeV9_]E0T0Me;_6Y/.)_NRMdg:3NV3>^==??1UV7Z]3e,OW1R;+17H:^=X341G,H
3dPS31)D@U.0)F]GR2N/Of@MUe5Sg#WG;3E9U2Q0D=P@G4J.:2)P=7<10?6DgLM/
#]dF>Fa9:?(:R:cWa#>I6=,COg?<0MXL9F);MT?,8&R_cd9.LK?R.bSVTgUUcSgT
65a1RTV;)P>_gN0W;SZ^DJCXBe_CB0a1_\AHg^N5360>aS.>9L7IT)6Q?61Z[O#c
Na#[RY]S,=EO]/[.,>W9_Zc#e2d7=eU46O(/TKdbLecZR;Da;^8YG]QE9PA#/=/O
OSUQS0X].:,7K))71S\f(TK67]<MeNV2.=19?C]=YaOEDYXPg;R+D&NOM>^dg,3K
F3UaVV8J_B/b-J46\Ic8=IGJW(/<;F)FI>\,MEDZ@dWX:I^Q8b+\/\TMBH)+WJ)d
0=8bF.-/R3AA/#R2]5XR#Vb?5Z68a66eQ/4L(R.R@KTR9Q#D2U:[-S=A56e:];&R
)P)a3ZY#DK.0G.6OY-R^Z=^MUU=PHPJ:NWC^#J,OMUbH^R,:L5b).;.837H3?.5E
)B(KW=]Y+2+1Z#OLBZUL]TD#<\.b9VbcU38[&)Q><B0:._TKc)-BO9B6Fa8_=NFJ
LQJE1bU0L8AJ@/.S(S;)(=15&8L9(:d[:1S5<IZ-,@,g\O6c/&>U-EGI0H>IBC33
eD_C58IZBM,8MN47:Y9a4^(d]ZIPV;U^La3U]Q#@5+[M5FAFS/+T(A:3g9eDRNBP
.1Tg^,:8G_aUZY#b2UR#dUWDQfMe4/L;)@2X;GO28QX:#HI_dZ^SbIa>eIRI\DGW
:0Ib8;]bWA:]=X(&aGJUGVUUMAY8/_:[O,7G+7Z7TX7Y=B8+0?SEZ&&^^3cBKU1H
B&]dQgMSe7C]a#d[OSdSd]AKP)X/EC1)_6NbB][O^]6K1NgCGV#d&BcH23b9T=eX
+-d=1V?K72#M,9&9)&THb2F4J;\ZEDRN^)UB+?Wc3;[6dCS1<A#0Kf,a4U^.G@@:
ePe^D>QV9c3A)UbCbbb&,eIU>1<75E?=GEUDFF,X>.c1Z5NJ#(c-cX-_LAfg,FZA
6DXfA]>#7gRe&Y::cf]]Qa7D[)61O?(552Tf3/)f?W5.,M3]VC@C@)=CQI7UL,C&
]aY2T71eF-22AWHU7)R[a1:;7;Q#:9#VOPM8:#QMSM8beYDb88HIHbN++<IJNdEg
M:H)Dd6E;:eINE1DCZ0)8Ba@YJ(<+IO\7N+F2H,TNLNBEKIMg^Reg/(2P6R4<:Of
HKY=U5:.4Qc26a:/:4M];?C1\:#_#:@3>Y>H2H9SE>?:L9+I2QKA)a=bbEQGIS:W
f3Z&Pa0:9;eE2E.7-McN-FVaZO3Yc#F8FC77U3;Zc-;?cQ.R&Q;J0-I)56V00c_>
XJ/Qg-gV6N-g[10=?KYJ/(a_8+gaDX.5;88W9,SI+J7RJUTCbJ+,2<_P\X3ec?df
EF7)GKMSK1NN4]5(4)(Wg@3TTGHQF1OD>S#HKYaQ89=/-@L,d278LQb^+\5=SWWe
g.U9E59.gX4f.;;SFPXWFg&S?])C2>f5.RC46W0:R(4]9O+/FG^(S\V[6G0)EK(K
+NRg7UZ/Q4>#a?d[=8Kbc=K(P5;C=5(Pbb[0OXDFd6XOH9a6WX\PSUXe-[b/HI/^
@<J4Qe2C,\>F:^PWWdJDEYM-0)+9UZN5dGb0QU#2#P>EQb,,E,F0H/PX=f+f04,g
5.40]WK@eW;aDKb4+V+dc0-VF/7OV>=?F9S4@GJG?FPGI(>c?-AK7,54:;A=_4H0
5P<,#EKRUJTGJB2^@?(=(R^TOG5@M^Y)8U=?7.0>dVePS^Wb/K&,+65U]NP^-1Q3
AF>eNL[d5MG3a4VZM(=YD06E07W\G(),EX(E_0J84Z[GbCgWM^c>]FS)6KEFR+0E
HVJ+[-QDDP04gFC8/62e]f8Y&8ZRaY9\_cF7\)\2Vd,:(aNXg<N7e+]??P/K]##@
87])@g[DK>E.&XUGbCNGCgMMR/&-L_RNYd,E(H++6NRS>H2^POE6Y^F#Vb[0#FTY
MSPR(S98N0)D9Z9-7gQ+5HgP1CDH\]=5PGOR,5Qc[3?/b?FfVB+M0OgE?(9-,_b.
\]YAB\H5d6D;bG8]F4DM,d@_TSQ2.I=IW_XP57KEVOT;d+1QCd;ZNS5eR4aG6@fU
ULIa684aB_)H.GWUZ^KQJUgX6&4/VHOgKUgUX+f]7/;(Yg^g1S2BU64gb3O54[-(
/9b[;TLPFWdZWIW)M059S\O\^BF8Y;g+/;;0:6T@]UAMD5Yd<LCMbaU+<7+.543V
Y,d.R\?3c?KH_V0.0Te^E;d-Y5/88TUdM5739U&/c>M9_W:/.&2SO9D]<12?YKeF
(B;^^gC1BG./7^^69;GO2a+I\)CX&f74JGH0/J-D/<6fb,M&P[=#RXFf@=[4&Cb0
JP]2XQgJQ<],<8XD?8\RI4\3@=?)gb)S7JFgb2eLUdQ8eS@XB<f>_\2-@(A1CZgC
BDG3^<g^e-6Z5+.BJ_9_(T\+>SI.I=b765;faccfY4L7dWc,Y<#B,GbNV:O+([RG
ZP,1dBeIC0#-4a;,-)(]gJfIg0c2&7KM]J7CU5e]6G1I<g[D-ZTUgF@A@0#aC-=b
0+9OLPOIX?QUW\YOHd]Ef+]aSA31[APdYIP[IIW+63b4WV0E,IY4dIf3a>OG+,7Q
V[Zg4d(()ZACY?X(KDO=.G+LI).EP:KBCA<DXN/VZe\<eC2A#dBFK<e,_]]2#P9,
49QbcT11_>.eC/-F5HEE)FR^5.cGN&<QGg-&U3FTR8TgIDN[P0(PH>)_Jd&8[(FC
2H7S4.82Z>F2(I3N&FbQWD1)+I&?C\d<QH5U,:<YN.cM<P@UP=JMI(PIF&FE;@Lc
C79dF#R_C]8;L&,L?M_IIX&/G]E39U#g)e(UJ4_I=-cgT/]-WP-5)]6ZQZ3K5._N
QIfS:9eX]ODST-c,-IRF^eYU]Ja0(3]aXH&[]-9EFYfG2ee3[^#BNZ,aW;J0FIUc
aI&/BZRT50(A5bCd4b\B1A8F:N030B,03R0d+EFM&X?41+G=#aM)#D^#;+b<\aRE
CNIF(&UJ4[ZAOQHI<SMd;P4FL-##7D[,JJ[Q9X2INGTVLJ1dZ+J\_-8,:P[BP#d>
?(H--0VSLOR91ZIFRRWa[I.WXUN3g_?]a4@bV<4K@_GRff<>+TcV<#[K=<Ab9e3;
4V:fZ\:d5VBIdIg3;&[Z1X7Og&YgJ<B-N>98=da(B[94U]8AHEA/4W<[N3T@WOB;
IF5[^<&R:PUE]?R>K?N/aAH5MOe_M=d&f^()/KM(6#K,GKRH6>RY:-/=Z]-7S:H&
67U8U;3N4b5=VEc(\/Z_b+^K+R,PdQg_&CZD@\CC@0+>/SOHOJ)d(6ROe?/8:\0R
@P1T,];BNSA41=DP^)?\d)_8I,Y\+F1<125d1RegZ/X8QZLV7;7T^PH;M4=[CFPV
-H[g_#RGc46_WVBbSQF-(XR7G-cU355e^.RVLdUAH=_#HK7JAdFabMTcT)a-dV9?
e0b?d6G457Ja<e.][_8bIJ:HCX;.3.LB]c.\FONe^]<GN-#NU=E\e+?OS9;V4LZS
H-/cf07,W5UO26_JZS]-cWA:\eZe9\a2YOZ0)Q,W?PC77/e4cE2>LT#GVP,P:gb8
CR\]S@<BR0PTAY8d(aM;6LT=,DD#GU03L<4T]H+;Z7G;^)FXceV@5\UQJ>4cE.61
0NUfbZ0#UQ/@LGHBEIM^-G6:O;I,F/[b;e=LXG6+bc2H1B/7H@_@ELB0-PS8Q&A&
_W8aDCJ&<1,MW0?6<]3(<[CC+R87LHG_L)MR8T4?RJ\3C</6Wga_KD1bb@9GH:H>
c9U\@Q/:16);Z3P:E5-M/<F_dWSO90T\>3gF47PbaB84K:,eY=\c>9^AeR,YdGb\
_+F\21\e</>4:VFJ8VHeHV,]J_a0]PB:2>)@&]7-)1PUabTG@?3HB]TaCFHJW@OF
>+5&^^da[D\9WQT.YNT4^BU#>O/66d0a&5&^&DC=A:b@<NUE8,#)<\I)[=Rd18H2
[8JQ]?g9,HO\CBT6UM]YYc=ED1IB9Tg3(?LM4g5X9\N8HK_#2IE.YaNDI<,:QPT4
0[2V@UMFd&N&)O9^(^TQaK..YgM8a6]+bP3^GOC(Ja,bZDE-f]dBJ.>^^#?C<4Gd
1C3X-g?5+.Q<4DI0L1S([+)>#.U\5LB3Ua;]Db0_&ECZ^Cc;Q8GfZ5d6#PfXWFE/
L-gXGbJ\gMBAc=Q#5b3A1CRE(G6620DHQT=@QJ)_/Q^:dN\WJ(RP-UDK^[L>)VO2
[/Y6@^],>QFN;,NXGQ&WfGGR)KCRRM2WL=D9\ceaD(5XD,BZ=\4Fe[X&YLW1D]c.
FeJE<^V>WXI>[HUYFS(&<=H7,98><HQ7OgGQIV67d3]@JXD>Be;I].\)&;=a;XW4
V8TEU0XORMRUWLCU_#EHX4QMQ[,]U4>Hec^Q]/G<Z&1PL;P2D(]<66KI?S3L,;-a
QaN#D8\A)9a3RF8ST52f>_CRC(^L2>Bf>K^:gD<eB+I<1A-)aL2(gEbC9P/(COU=
BI5Q-OA/:@f.=HOJ^(Q)-(#Y>&/XE#^a3:V,BM]47d+,-?4[12KN/6[\I4JSUEL-
?Y80J8+/@IGbT?aS9FG7.W0c2Zb=Og8TR\]N+\5[<?Q6=aPV=8^)L^Q3)/8SY&3;
K+^NJHNDJB:-GO:4-AH;_;-eI2R)=#R:,A7X-F2FLQO0T&.U.e4P(G2^FeO7IXJ&
(-#AR#Ec^NJf#N0/.HJ.&\GS/+P-7a;W=.C51JMaVO46@g15ca0b><CVJf-5/W=e
:YVAe/c@6)c<3\4f-O8,Y5RfVg@D.LGK5OUZFW_85[&TeQ2ABF/dK?c)M-WY)97J
1^R8-d[T0cGW(R_I\@C;((S7JEZ51?A;:Q@(2dXK.ZaU\TWPW/\+dbH8@HMPY8JN
C&g?Yc6=U?-;NaFa/Vb)T-Z]M:BDcMTSB:S,-LYTY.NOJg9IHM_B&QT4D/>U#7:C
7:WM__.)?g10Yg@Y^g1)C,Y]KdT=LWV5TSgOgfOHdJIAd.YB_,f);JJU4a\)_XT.
+O^;C>3@J_LI#96X_H3Pa<2f53N7Q#X<-/a_2;K^Q_B@BIOAU-WW-E9EWXP93bDH
MB4P42VT/@9ZG8N5?2JeTfD=)AW^QH5XU.2=V@9I\:\c+5N;S0#<0+YYE^:/9YE5
VaaAD[:I#[I1OS<S>5SW:dAbeTdaOb2KU0E4aVU;FXMdEfLMRJLTJ#7SWWL(HZeS
TOf<F67WG(g53VHSXQ:86WXJUV:CEG.3._BU4AMWTZX+e#JN7PHef7\^OI^+K,GW
g>g_6,65V7H1(4NCUaK_19&Ue6EPgZOO,P4WFVR=b,Z&IJ;aJ5/.XEdXK.LfW5Y+
ERU4+JH;8G)K)L\+Q&9N^HK_^Q3F.HJgacNP<0FXL?\T:\7WI[9NADO?>8IK&:/d
3,&V(ScJ,P@#)bKLHEF^]G-&_FUW3E0NLd76[GCYb1^/[><LX;dZ5Q+ID2WaCRX>
8e1OM\f>MWG4_^:1/XI]0=4^[=DAVNaF053g;69X[aU@e4T-ab<L>AQ;B6JcgP2T
D#<@P_^^>@_P6A)5Z]^Z1;A^c8.F/E==#-N?+6cH5bMTUg&67,PUYLH5fIDHQE/R
ZYK.^^H>PeA4L5aX9>#MQ>GT[Md:UVFF@HW]N>OS_M#Y6Nd]CDEAQLSec3K7>f&;
31^:E+O0DNf4eJWDF4)YYQ8[4bL#cD+YHaHB2:+,^\G(;MXK2+]^3c_LX9A;MU:8
]ae=^ZUGKU#0WRF.V&N\+UL6PRV#+bI7,J7/E;(=eT^DVG\UT#dNJX>H=C#MP\60
U+J96/8bE-.S@ISVPb-X&&S:AJXG5XG68LPAHNNS[U1gLcY(S;A7?)OJ,0]#c0:Z
QTNY(Y+91f7@?=\DZQ#08:R3D;gDAX+L>0CMbS0@WUFS)Xbdc6=\)-e?9QQ4&+>d
SLeS<F?\b1LA6TccB?W,UPTE[JNgbQN]BPd__;:JbEAa0&=b_QD(,eNTH?OWS:]a
C?aNHD&.Y+<_B<1\5O[/8K31Z[aT(>#/@/J_9/5M8^BHI_+YA]SG+YTg]egV&NV^
H_BE-R3NNf0?D>LY]KT7FP2@1fZEB9+@fX4TEX5gCIcM8[IA?ZN#P]/I;g\&Q5)2
9ER>&U4_AeM.9YG?aZC._;0-f_^]6O6+]8@.3KW3:BPK\(<K;N7@fZ#74=X2#UUD
3?FH^S,]aMV_EKMH_^PXdL@OW9]-_^BYNYUZ7C]f\a=@6-=T76DTg1aNWF(\=dP^
8KBg]R^Fe9b)-I/_afH1d2c9f^\c6dZgg>V.UR8S)gK+-/F/<eKIW(FWF^VcNeW@
1&2:W3BT^cZ^1+Id8^[^f9BA9R=eRJdW4f134Af+1#RYe_f9W2?AdcYK)FJ8[,c#
F7.G=0R=GG0W.-IWC^9UL]PM;.YU/MVe;NEO7\SMSZZUGfb_[)WBI:&(7N#>EdWa
]VCP=@0J(MNIH#)a4NabOULGQJMS3,_YJXM<BPVW(^>VK_S&-Neg<_K&F5Nc3?b3
6E@4@L+U,>P2&P8TJXG#C6\A9fH8:GKOI9U=cD8bV_fdX=WTWIG8b-FK?<1g<T7f
IfFCEX9VM7_+H=8=OTb)aJ&EZ-#CMaeR4d>C(U_3ESQADG97C,V=gd#.S=Q:R<bF
LJU33dT2LHA>H30;MXef3(_0@8ecg-eBg[G3-RR1]=fA1N;Va=#?J(25[M1N4:LD
OgFAXab_MT6gf)66<Z?E7]-gN?#)U=73G5)6CJeN\4VY#5JeO]?OEMW;X:UC7RG^
&2>XdSG>Ycf9ggVN+bK92OG:62@00f#8)S2]BS^_MMM\:@@52<eQ^UKa5WBZ5Y:V
eBgFNX+D.Z(T9CT;/4OCZVJ,\3/#LW8240==DS-[W1MV;gBKRb/F43?>]A+bdNZ@
W::cXPcI3O]?IW_@3TcH[L>,RRE5/_,VPOXEU)NZ_O5C4<-7NSDC]B)NS)fdS;3d
#\?KR3^?O6?#g_BY_MX+NAV2)g5.=OYA@3e_(:-IMF?FbCB>6c7P8B#2G+@ER#b;
]99ZCTR,b<]g<b2a72]J4G\)F0=>-NVG^cNd4\7XY]bR<MP=>M=K\b]]>c5XUc9\
?Q_C>&15dH@[+F4U60[QASg5U:LEHa2+8;9LSKI7^],686-H1556T@@2L5Dc#25F
\DZ_SDg4eN2^&)2>\POW&>:cHbZN2M\OIW\LY](1WDcMCBd4KQH_HL+G<K8G5ODZ
I=]&8)=0KdK.[:#+b:J^1e<<A;Q3#][2EQ[VL8?ES5d.T.?\be2S5SW(>MEXTD.A
Gg)BGSU]&_VJX(Ab(:))R<:56/fF0g6(a2OcFABA=L(3-<SY?J_)Z)7aabLCOaV4
S>DRG:KUQ(.BRdSTM=N=W1)bO9].R2V5I#<[dOS_(RR=:Y,d3eG:^70Z^P]fPUg3
[X2F5T=AQ)X3UaX&@/_[J)<&\>JSCa4[A^WW65,199@]-3TfF;>c>-JNaRT.g[1F
,#cbN<5TS2(G=YfE2MS.,[7M8.c7\O?a?ff)aVX(^c):L3XdH71f;7:)LVW=GVWg
P@_6G=KOQ/T9;/7E.=L[L4,UQbDGa4W^^V9fRVc:C?9@1=&Y,g]d46>=AGY[fVFF
VYTbS<T/?TcX2/+P.2/2NR#;))R;cJbDFB[@&Nf@g-U[N>]O?\]4(:bd#3/f&MI?
6@;SW545]c^_)-(K/6J>.K;/#DX>g@fb46Q_)P&HV5aZ0<+T24TC8&M=F,;@@;)g
WS)2MFgeF;JCc30:H4/GKDeeMZRR<TITdMLZbHJ_A<_^#E#IQB]E1;58A>ecgV.A
IKRaH,Q^LHNRO>T(]&FWN>+\[[T<OAcHB[;?P1C8N>T&XRK,C.aHRSc=R3@::b90
T8W23G6;I\VD=d9LH6D2BM<Q93SNA/=f\,W8b)#70.R/b#]DbD?IADBe/KZd86IU
a_X#<G<1M-QTK;I@MY>5IQ9\PQJ#7H_)53C4Qg]T@=XX\,J+e^-de^feX?D1[R-S
[&><6R86PD.U,-^M,BE-E8A)J7-<9?U5&b@W\Mg?YEM0,W7_f703]Hb94Q3U>C([
6eVL#A>TT/a.P.,]M2SFO?,IL(26,F_Fc)E/0B;f)@d\UI0KdW;S&)cgRV.HJYCL
0:N)X8XN::Q9]EM+/UE>R2FL4QRP+PC+aBe#JO3N&CGD:@===f<.D0d./&FF]BHK
==\SVH+fF#@K&A8+K9FB[_XUd:7URV@1(;A&WN>9[]Q>8#BdZ/E2A3VS+??7+Yeg
gQZ.c]8:T@6U+0\(#J\/^M#LAeGQ.V=SJ:Eg<3_>J3&2M]41Z,b@[cYbN=f6#9]Z
U;.[I#a)?&HQDB/(T#bH6>gdbE?;L//\J=RQ1;,M@Ub9CZY=]QPKJK,[S#gcJb.S
gI^VM:8+^5/7#O<)+d)aP26ae3g>[,c]@G)>1XI^F)H9ZWY89I#069HG^TK8fDL:
VEC,WDgS-X_/OX?RAD40XM)2c4KMVXFf=AIO_>WLB4KBET=^\:<g_cfM3=g2+Jgb
H^QN=DRH2J(+FD;X)L_TcT2?D\dIgDS=>0JS5\Pg1VNOR^eR@,3]RPD<6Z]FVIGB
Y+O05UCJaE\1P0eW1\.P.?.I)G2A(M[K>3ZCWfI?,A&dQWGeY]<8b0PC4DQPM>AH
4OLYX(R[eaY=NB2-cHB=K75-<L1MEb0@aEKY;fQ1W8_?/VABYZ(:N2OI@NVDF]??
QQ@T&G\4=559/D?e_0I#7b9:/9+7W-]886JTL)6N,<=?0<@5/SaH(ZEPY,)eV+0-
[dM=Hg6QcPMMV=6c51(\S#7YGQ#A#\DY9_dY6\:Y.0IJdO:C##U62(4g(6=;A_d?
^<Q+/HFf(:?M@-2A;Kg7bFe#>K/dX\/-&f(V4/f?aP+Q3Y7MKfK:d_:I/YC8:[Y/
9X5-1[c,IXZ=a][C0_/3LC=ARFCA_X[5Lb@ab2W1=X2a3I,0EfgS/.>S3DcDG4OF
d(g9C=dZS@#d^X6WKg+@U^=[,=0+N12;1.R66(M[\(.\6e?dA2X0g<Xb5]&U4HGS
YPOR9___ZF\c>\:da7SOFeAP.2U\a9\?ULS=?P\ZK+3),K?C8/V2QfJY94EJe[@;
XHGWC0WH6@S_gL))>9ZM:H&U^[O34?Z@<]a;(XQAJd1gTVKCJW[97WTggdA=gF.F
cB[JP;6ZJIEECRWWc@QS]R,#;22.]5[eKL/O&ZL99#?UHICf]>Wf(Q)Y(Z<XE)Ea
;b^5AdD(?&Q8R0YKP4Mb,]S5eaYgadgY<2H9P#dQGV/WZQ#b^Ka1;BL#\O8)HQ(Y
c:VJ[9J:gd=KdC9L\&2GEN;g5?8;;]<SCI:S)E\WR35VR@E^9#CS)?RBPUKc^[7V
a-c3ZD4c#Af3)@8YT-(&&M[4^bg@>#WONB3O4#QHe2;S6)6TKU<)dE4K&4/gE9P4
(bb))?HMQEYd[b/T/b?=P5V_QLQSVN.Vd7=?&d5fSMI?ge22,[1EZF-L2<E@OZ4G
W/D)V[S4=_0e+G75-e9\.A)20(2[VQYD(g<bfUYWX7JU&20HagCdI5F[FGP)a+b2
B/WP_#NdK6L<>\7^R9[JEB.MgdV>MD4I+MK00d+-Sf6\.-^UDI@)eIG7A:g-0/^L
[,+BV8\BR)RL#>O.\,dX_U6B8aC2W2.23&>+D?PW)&+HTV2V1bHd^3W40IVF\G2S
B.^1E8Af4B@>>P[cd^H#Z]4fE-4PVEb5M+/W+IaKbB1]8A8bV_\\]B<#AaEWe=.F
BUG.b]_OeAa+-e01WF@Q(B2((3dB#C4A4N=/+C<WEN+O;A&,^VACL5;2^_0S>[IS
,[#SV6GS-\_2EfKW^Q,a4V;V)D4&Z<?/eHZS9I?U29]31I(^(3_c<H&\a^9BbD])
9K6>W(=A4^3e-MW&;YeKL2-9HdgA;\[I2^S3=R]A[c#KH@#/;A3b[gBF^.OK^UW8
.C5]OU5P:bgV-]_=(KbBQ8VdJEEU>fQD]>e8;\?Y#E>8K9@Eb-BW//,-afHI]Z74
1:-(QI,YGf#489JeL.3P)eFYdQde&@<PBdKTX2&JM=FcN<S844/0QFLHe.H>R<N:
)<0Gb2UQgDZ97(Z#MRL,FLL=37[T0>)PE5HcNX5QW?HSga_/]fH(\RJG,>KfF0:3
3>AS#>[20Tg]OOX#d,@QU4IP[/=2]M>WP^8<OM1SZ#Ce54ZF8+c56QEcb2G<289:
P?)X9?V2(@&]RGAW5c=dg0e4:bf[\N[0U4#;[GKEP2bQ1.CW:0F^YP2?d/;<FFF#
.bV3)P3Zd_8V@)WNcB-EE<#0[=OPLT0&e0/;Ea^2ZSb9].?TXeRVS^_;CZUU.1SU
W_#2>F9Jc\eW0<Ua2Y+e]#a=^Y(->K&f0GPGJ8YJ\[W_.]2KAE_eUOFP?NY:RI^H
GF5.a?6.<TMD<<=&^A&:81<MBf<E?.5MHe8INJA0Nc\b2\5[[(OOc_1c81XTLA^&
=_ebGRD1]f/]^Y@&]S&MC.:J=[/4;+6B&S\Z[<;8-\[B1b^P>.R-_-gB+H+I+9b5
>U=#[#+B^Z)T8.6E#71+XOdg4:X7H;:?6(D-?b0]ObE?VO@+:A?.N1Ag\O3L460(
bYS/H#C7R67/J\QYHbTH>SVH==C\ML?TA_I)53BD&U[Nb^R)1JED^F3\7UPB4HE?
.RcXS&[4;24]OX=Cgb7,aVc9ZWW\2O^;^5MKc>9:<<56.-@_&a;U[eP)5U=P?<Rb
DT=&43Y#YW&]2#C+#]XJ?Y6FNd<dW-69RG]\H;(PL#f1S-I9\4&HYGadHMVEIbHE
\X^:aBP.b@)T<X8GZQWc)41]K_Z/VD.Y0@d56[Eb\7UI2E>Eg/a&f?^gd-]5\#NA
<[K]dN\aQOQ3e@9;Y_?1.aeMWE&S0M,.I7@HXaL&7SG=[/F\gUIBFJ:cc]P/W1?:
D_5;10\]#MEQ-7P(WF;I[JX9FQJ7=P[I5B:f\GUS4FHDWeJ55A5a@_?RB22<-XD_
#NcJ<CB4Q&ZE#e^34dC.PGef0>-CcIS9K^<d<R.IZb5DPSF(_fP(?^6;69&aO7f>
?)S;;SXNOGH]X9gdKOY/ScN#W0N^EP,5_/7X=66X\b:/]U[8S[C83-/bd1\:2+2Y
B]8X;CBCI]32^I?V1E,ZA:>KLZIQTA?eM>/(8=[U@32YL2Hgd65c]ACgG)?01a9K
G)6/gQX5M)cZXggFO<&L?9]7,_Pc^M/26M_MW)/JPWDJ:&d2JG.b5M]2-7A;M)>f
OU(.]&>Xb3^1QEU4T.Bd6_-L3OLVDLU1BI/]N.M.4HU7+6TBT#9?/?L_RbC@0EHM
>&&M14^(A.K<KEC8b+CgbLE)3Vdg?@BEXGY]3Ga7gZ_FAI</8g@/,47_4R(bg44\
QdXgFVU.f8PD3NP)EGN_K;3UBXX0Ce+H;K9CK59XcIfgY/WJaEU4OWZ2(Jec&MXZ
gC8G3fCI@M[DWE[6Z??cVCP0c,#1\Sa1GYA:SfDVC[\4\MdU>:FC91OBb//T2RRD
1cfFMb+8E:?:.X]PP9PJ/\J9UY<J,=HN69(MI5T;>#bVLS/(7X]9abe1L(-#)4:4
ISNgL\]9M=.C9FDYL[6)F,1T&;HHJM:4+Tb+Z4bB?I6KcS_<g4T4-fNaK]=Y/=\9
K-FEe?X\N@QI4DZEPW>;6^SP:_M382e3_3&VX8M#.e@W<a[1V^c(64fC6dG\SRLB
FC;H<P#&:D2.43V//d4CYDaD+JP16E^^EDJUb,-MR/e.H5RIA5KGJXN-T5V&Tbf=
Z^Q-aDZQV-K^5G6g-:7GO4A8D)DY^-4>)[?5)@:GgSHLdZ2Ff8J@PR)8>gZQ^)\3
MGGOQ@0ME/8;:#(_Y,HC@RCLaIPe;_0R@SM]Nc^\U1X>FN;CRR^Ha,g+]JVPYJ>,
M:]@5^JJ^[>M^6H.Z_&c3A4ZD1XG+;T?1^PN8/&FM8EKHR=9.Y8?HcHQ\E?YMYL_
8Q>D\HBdc(<RBdB=?PUQ\WH5EEA4YU-:^0#1DOW]:4T</J3Xb2;\A4#9D^6gc7MN
#Q29IRCa54cAce&,=PfV<GH8_-5B8BOO]@KAS4.GbI.PI(N47C-#UbTdY4&=?2?8
M+PH^=A41b(Rg)e59FHOJ7#Va&HZgV)LTM=0G;d6O/YKFC(6MRHYXNDLYEZ.JcSH
2N@F\7[P8>c\=U>_/MP0MU\<OgX3&70(O+->+]J(d:_RDO>@6<T5G^eQ:dP5d[[W
QAZ+=Q911=\?ag_aJHeG76N93#)d]S(#5G;YEg#^06f-V?DC6dd6Fc.55.2QJQ6,
b1D8<P6VS1eS4=IE?>=EPe/3C+]8GPH2A8?]/,?T_=DV_(;<H@e[(cHD@&<fP/<I
6BL_bR==X./-f[4U:F#=2IT3ER(A:;H5d7JECOL1f3([]PXCIC8KL195(K5[ge1U
F(UWV<Y#?HB:EAV>FWNW)(+B.H]:M>fC0BNDX.cLQHa.=d6P/YG,-@+>+L2XR9[f
f-dY=Ac0_;ZBbJSWeE])8,I5AcWAfX.X7DK@NXaaXce[_WQENK#/#@D=CGCQM9ba
M[I21BKL_+,+@]4a,dU0QA/ANAg0\@AFQ9)@S8.&,2cTW6-Q\:)CJ<,Lc/O-@SY1
O\M\G0>?\8VR]88,f(>c<[98e=ZLZ;Q1;5g]0Ud-)T^>/6/RD:_NG^TXaV?3#4ZY
b3F)((54R5JIaM7dNEH2<Q@/N]#6Y/1SJ)B[<^BgcUG1S&R1BM3+H,@G.VP9/b.a
S7RbTP)^:NU,QaQ@EZ\eLGVC?-_CLUL;XBX0VD5_&fa-9WD92D;OL3A,S):8+<UH
.aa)44GB]PS(\QVCM&0@?/<7ScY9MJ4@NUL+.a-==JT_.D-[^Z]S9aYeRSFH/KI)
0+_3GG]J1Z#]aF:O7Eef/N>\IeM3Pg3)#a:D/A[OQ-,=)Y-6LJIX]HR;T?W8D4T^
eS.5Z8TRC/F1)R&AK7LUbIXf^3B[S?]=Q^R@&JUK/OI\/E@;f_b?(D+NbCO#BX=a
L@>;a@^a-NOCMJBbcBV8KHB\KB@[MbK7PC@XMJG+7)B?R_Y;26G=>_6KV8(T]Hf.
d5X1]SWW:F65NX<=c[4,XgSVGAEe>YT?74eSG5f&^<.;7/a++@>?(VUFW(VXR_@L
-.G]\,OEMREb;[W.UFE,:#(+9SFcTHX-N.]bLR6gYE[@8JUe+MV>I=C_Lb>DM=ZF
F;?MHR[3K+M23-XW3N\9LAWEE-X#\8Qd>CY\YCb##3ccMOd26CPg<0::\:_39bV@
V+\2>3UHXSTf&Y:O8ZP=50)UXDOA)GGFB-f/XH)5@BRMMX@KdO^.#,]K/O0IP4J4
+9RP>59cC9^dTJ(I<989BBX>VZUDecM?DBV,DR8=00EM9dSAZNRUa/E-[V9E0bF5
)2[bZF8#/PJNHFB^>;c[RPf:9V&K?fcdQgI/6X-8@dPQ@7S]GE>#:BC_A5?M198/
>:&a5^L<Y.EW5aO5ZMe4e/6e.#f;(N;PC\:#-J#XL@[;9W+3SA9?WOPQ@gPU^E2X
dYV@EOC#&]gX-BG/3]g;IMe6ebXMXR;+?,#,?Sf)^IGLJRe#c)W.\SX=IQg&fMB7
>Lga(gL03gB.DPE1<6Q71bTP7B\9@FUEf>8QcT:U.+XX-gH9AJA.4\a)WOO56.SU
Zc3BI(^@OfZX[V6&_?cKLUAg_N(S2?V7a,-_>2:a(aD<IBWVPe:-JUca3b,BReK6
TC6eWP.E2WOSag2b5[cQ9;68K:LSQT\g3,/IfgED)?@IR7V8>S&6#D/ZD0G/8K7X
b^_4eXA&EPfG.CZHS?gO9;P[G7G:dI21S.a@ba?U(eI[W^[+M23406f33X]DXWG\
A4TOPDUZMW]\+[K;LKc\(=[+7c-5GC@b+Hd:;\(Q[H\+J?;35^=G^[EO#H-:D0=_
,4dF9X\1aQ(N]I)b9c[Y8T,Y:NO9U4^_.KPg)5(KMFM_5=(=76?RCL=Mcd3_)RRG
6Hbb#Y.YfL0c@IdXf#_b>C;J1RVPMfe/U<]?[26X45.K@:Wb+G7e)4V=BC<1ePV_
)GfcKHG+MN5C:X3e8#2)2g)Ff/8VC63DK,B1gNH]T>/56YU(E[)?[a7QDf>Z)b.B
6)_1fU1,Z5\L+0KVY#I<64AYJWX2SL4ef)\CG,15HL(:9bPI>eM3KG^,0-)VU1KT
ZO[5_d+\b5E5=@L7-R0?b.WP>)2\Y/1;^dU;4e5Y)P>d<PAE851[bR]12F-&[4DX
dH2BW2YC3c-^+UME4bNOHCCGcLG5:(F5_8>aF\C&L=gb?-4A6d.H:/K==5NE@7(M
@fJ<ARLeB=\U5YRf)<KdaIRL@K+<\U:MDM1-Z<,_+?F<]R?>\6.V0#fK>^)9D02g
Q=.]7S06\7H.9F4Re023[_Z7@Ea3(&]f@ac_H]YYeBHD7:PdFJY+LP8:GV]#S,FR
Yb6b8(7P:>-SS:C;<0[e3a8\/ZBV;I8H@(^-c8&U@O-M&/;b5@eI=A9K29R1DCJ[
9;HZT=;CTKe/KZ2#W7D1KIBZS_\e/XW,@4.APKJaARb0?3C6T=:_dY[P+d:-a1Tb
PS^cg_-QL6IY6/_RW<Sa[f&);AfU]30G>/f1@>OPF0ZMf--+4A(I]QBNO[].6;.<
CYHf@U/aKfF>GM<BQ9E5;,#&LeDSZ?&eZXUC/^SRF<1#;;BP=-(B2LC<-TU\1L9e
]L6Q,4]EM<dP_\O?Q==gfg:dA\A7P:Q:#/S2F]6V(3W+NX,Fc+#U[P5,eAaE1R8Z
.O^2_<:X#SKC?=G65^JDDM681,0./ad^00d+AbVTGV@8J2#;V2NV/>NEdF47d@E,
WW&5720N]==PS_S,6YMO6.YX>D[N-R23,Ag.eL.VA[f1;X,:T+Q1PUB@CgG3UQ[)
@16Yg8?^[dZTQCT_&,6-0PJVNF?=]G8bU9K16fdVGJK\T[W^=TF9XJFd,P_;WKf)
TOL#=8B2cDU6BFRfVV5HC8edI87aYBeAYe:.f0e9[E&dQQYK0Q2KH#:[#[)_@KX6
[U^eSXR1B7U\W.a/39c^CQ0cEJ<Q#gE]/_8LdVV<F>(V0R=:/57d/&<Fa^>CW.9e
B&^1+BMZ#&-RL:L.S96VCTPL.fDeg>gASCB8WUJ3>F/3:P.HB;\c&\<D62J3]?:W
^JE6NK1(1#b2;[X[D<T]EKP+U0cIB<_:G@/UeZ7B)KTR53EQd6XOYAA+N6S<CMYO
NB#59T2NAB\6fE#G2D#6HT2PYQa#eeKBGM9PC(I00f,9cfS#0ILE?T-I^;TC::H[
3,(/6/_#<M69>#B?Y[Z<bZ/=5\@C90[I>d_P)<U(P&_#R7F31E6OUB)T3&32Q@/?
gfUPN/<_TU::U[M76Bf:F=B1V-4Ff@AQ>_3_./KO\X<EaCVc8G4R]1S2eD;U3f]:
8B[(Z@+FJ6H55\RX#Ua8Q;Sg#GUKe>;+G//^:gPWfD&KBA_R#1P3L+I(I\[bE?P7
XGK0d.QL_-S)A]/_#9(Vd\.eZ(X8\YNYAB3006:f;66(<>1VB^f^(/cT,K:\M9dF
@=b2A^F^L4)f<WTO9aBd6#TX)-(d9BYMG7(+OU,2WY3)EeL=G2FU3fE2(F0KN35J
#dUBTIf;HCN\c(Jd\)+@S-[JB[6:EJLW@)F+IF3X6I/N[g2KD&];9/=<#2GBFEV<
)XD1:)4LT6^KBJ3<\2OCONUNWC@C#]SUF-\?3LfOS8I<D,71[c^cc:A\;4]IM[fK
J.CIKZAFEV/Ya?:MH/0aEfgT7cD64NDZH6\fHS/S;2d<LPB9=]3_&BdI^Cee61X<
3Pc)gPITT;67DOF&3HX0I=ZAN26O)T>08&,N]\9gB<e?a^0>N-7Vb&3JP3Nc/K6g
IDaQf,D::1U<R,^6:WLNgbCBO^fD1AD^a<0KR3#aS9EDaZY+6=8C<<_H6B^YJH2\
aQIa>3@X,-b,7<H,8,^J@Nc]]H=)[QU,0Z?BYB55>a[.2c8FD1c\cG[fBA<\]V3K
F,&,VKFWD.N&]B:?UR@X=AZKE=D)d]F)dXgeGZ->E]F)a[VB@=53-&.EBEB]X<.8
?cH6_B)B2d_>E+)JI\6Z8b_PD0?QL)6H2#IX39VOOF/J(:NN]-W7O8QfMbESJHEM
bX^&IL-6QQAED_?H2J(1<5UZRIPHZOL?>O^GZ7\CJV[A6/e#<U2>G/4GQ98TLO+?
AI@@:)\KagbJbSZFDb1MCNd&7VHRGa)EeO&KLSca/gZV&1=R\O=TD1P_g@/:@Ffd
1C\e&Q06-?MX@)NQfg12F8cE4HZ,ZY:/dV9B[QD@0?OfC3?/+1<P<&g+=(HGA2@(
ROJT>NQG)K[Y8C72U?gD^Q_N?Z[/?2Z6Q;GJF8bES<&\0I7E^N>JU;<bb=P5Qf9D
#HP6,?fg<QW5J(/0S5M+=KdfZ[#V=-O@#;2/EZBTQEYKMT5J(=V,Q#\D&U#_;DLY
QFBB;Q:,VW0[DO._fU6I\82^6=W[A6-;O&VBfF2>Fb3B>8)g#(cK&:?N@bFQRI27
9\)0b9d&/[38\<<A#BST65;()C(3XZ(I=>e=&.e6I6S9TId_S&)gPKRJ,/DHbeIU
W1V>dc1HWW_J+V)[cRK]MOCPd[L>J5:3gR6^10J5>RTE1;Z&:SaIH;I?P1WRV>,M
D1N;2FZ9H_._bd6EWa[=1<@9H?<a)La1TN)eLe\G2gJ#dS06?WF\.+e/<ED\8UbM
UPgDd69NW?1G7/=^\I0>Y,,+JDI\,)HGAP<\6-3-\e9bV7VdHCJ/T;Y:ZRNK2X:3
2[S#.;G5KNQeGNf8-Z4#32+WPX<GfK<\]]JV^8V20>;,:+<5X).EJTSO:GH<XaS3
Y7^W7_U@^9ac-Q#e3[@/fM=^[)\L/e;T^W<5R32F(K=9^(SbFg&E]7Q:EF)5W8WQ
3&;4)JVKUd#C>:SBU)FD-^bT;@?90()EBP9KBdV]3^f^@KVKW5<@_Gf73H9ZT2\(
@(9H<A>K>O7bAH\?g9C]>\#8NK](X\d-NG6NL,240OaRSb;OOY>V,>?2W6&VdH<:
bCM4F\T2.efDS045eW5/H,QN5(;P8L4.10=3R\R4bUGQ)ORI\HJ:C?QA1U34<Xb(
>W;^Z^X93[#Sb/:1IQQF;ON?YBX)^12L(cPYGA8c<#1,bdSVT(K_C/4ac]NbA<5;
D[387(C3Z^?93e<eU[Sb8>?=SGNeCDVc=g\f5&Q0cE\YRODUY+5[8T&:01&3Oee2
4=[Y3D6ZKR:T3=VH&W=bV1;P<</M]5;LgI&=W/Ja]VCQU+;1;11.GO(RK5OJDGN4
;ZbTca4?<Ha&-YM](TebCfTM512&]45K;cBVPDd+(\DS84OMR:M(#2UB5&9;,JW1
2,Z-652[&5<:L27/cc_1M.5VU+5H\3F>OY#+NMT)4cbHC^>V4O#OUL@5C])fPKC,
46D+\TBY]BQY3Q+J4Y1,CW6M]]@1WAC,#KaQ+,V\E>5Yg1T>7^PK0GK/Q/>XLV4^
@LRNcDC<)g^Y.G=4Lf7bQeB9KM&56BZY;W@WbK-XADd9\W3Y8/UfO?S@TaJ#PR3B
KFBQM70RZW2XF/dgB=JUafUeSV;T\UJJ[+bWYXf2D8?[0RW8;b\bBKV_@+;<A&RT
_R?F[+@#AFY\UF)W?\31J5RC15BKgg^/[7Ke&Zg/S#538.0<2;_GUYY\gS5LWZc0
4W3A[U9OYQ\VQ;((dT3F/7-d\[IZ^.,E96>8;ZbSP8b,,P/#C+d,JC45-,R30P9M
N2@@A60If^/0-N.M[6YaBTAfG,:cG2L=eJec;1FIVIG734PA^?=;-1FI_HgRO=90
XV#RVV^&QI09aZ-L[-4cRWa0,A89PUD<TTgBISJK<VI1]CTUFAAdHS^\AB<.Y\Yb
.D]+c/3@BbOaIIKU(PXIZV8YF4/3VaNY:3>RQ3B@LOZWUb=+]Nc757/DOUPZMN,I
+__(?@=S@FN)3^;-DL#H7NSW)I@Fc7BCW39,g]AZGZ(&J?>1+f4#S+e:K)gG^KJI
KW2#X=Q.WZ>5AN)a(MSYQI:22YDJNOA<,\&efcJVQQVRP1<Oaf2f(\^MQOHeLK\G
A#N_A^V[^707E>#H/Q.MY[KZ#cIVKR5EX3B,H4cJ724/8V0QEX<EY=Z&:6_X:-0a
U2eL]aWd),;aN7J1^;X&.490Af4;]#FHfC,_ACS[a7f>52#Ce/P6>6Of\Wf.Bf>.
ZB:(Y4H_4S3WEQP/P;S;>5&C)cRWf/O&<gDBW\ROO=3CLg>IKHF2H(F8<CZa)K?&
27fL2VggHF&,C1WV[cW)DH8KHM[7\1WG5M5BCZeDDU+US32AHK2:2eV_Wg(/_O1Q
R)#F&G(bb/X[SKS8CWZ&F&\F,5S@4<\PBMAg\Q\)bVJR^\ZA]#_8)+^]OXH)b\dE
KGL1CaBf^fNG.e\O?O\_F_^8,Z<Je[F^ZIga5F0[NA/\+&f-_LR;&W/cb3C#D/R_
RL4,TIaJG<89I<fV=TF62QT:T[AdHN0gU-.8C_M^I60,.9F+72I1Qg[(cP;9f2GX
(@D+NZJaYT7(5JTbQA=I1b7R_^#C4N+?(=f.^L6>KIA6#]E]I+#(cTU\WC-YS_\E
dB6D5IU,N+F7bK9e?0J.HS?<\E\YVE)7K;<2;4VMF&B4N3(7Z.P.4T?&A#W+F,VB
J:dS_U,fT&JFPG.Q1/<1@<<C;,<eU0B<@&]KW9eA?IX5)V2ZM4Q\D-M9#_bNI4b3
b6JMP)0^NGQ,fM<M.=f&KR:0[./N8LRR4&g17-9=aMd-c&/Q^5<+K/Z^JMb\BN_+
<@I4d7;IfIUSKH713g(Q:@SSJaA<MN0G)/Y3cZIN<<F2_JYb7IK[Ie?R=,RIT)80
NdHPM^Y>J>=2WAEXDM+F5RP/b3?2:>8)@/A/TDcgOOP7RXD7OH]QH:V(dbPf4XDW
UPXTfa_YDbG#AF8a=b2SGGXO?I>f+\WLMaD73ZM8=ZWKK5-b0=514/^:NfD\Ed-8
a-W40-ENCc,[1/_Q?[@]GV8<KN9O>0CU[e>+RQ,2.YPLXdYK6IKMBBB)YbTU[2[8
(fC.HZHAE\TbL+&(MI8>B?H/7+;DY1^0_b<M(^c54ad?6\.N.A.[-)7,^X.(1EN]
8T<VI6+Y18-2O^>9U2Cde,(/+0YE9f#?E&U6(Q30G#-,K&BQVX_QX42<BH,L2&de
B4a6,:bI</c^YUa3RH:?6a<GUGX+L<?0_(#@)AG:f21^X.62J4g;UV4WPdV>=Mfg
d.cHa28@<<^O7PHUeFe2\H40V]SYY_65[IedUY9d.Kb>TggJLV#d]].e5e\Q6K6d
2HMELJ514W7gg#;>;DMN98KYa4DW;fJg[E8N-4Db-/,Rg(L-_SK;-U+);b?&.\Z6
Q>Y[[<YDG2/YL^=?N3+S@eA^gL,,8STZaMFRPS]9-0NP]OIN06I[8:TT0G87<I.f
gK>g.JG4eIRBZZe?1X85N.MRB+H\;NY-A4]^:]XP.<&VK&abL_-CT#SMR_Q^RT+-
R^_+8C<;AB@Ldf.6E2B7B=)E]/&J\DY[5-VGgOHOMB0<<b6;JY,e:+V&=\G-R4Ce
[8+2,f?.<>LE7OfOJN9#&T^0:Y5UPcU(O\:MK.J/R@gTf/&MH&T5;Q.,K4c1MaZJ
1aHK8>ARc_O00<g-2<[,[?2/4FMM)Q8F44FPXTX.D\,bQ?55EUAQ/&VY;\@PO/AE
cEbgdY>Oc.<B/=FBbZ<<4LPa>CTGO_5eWDA2+T,#WdY#;6>L8ZK4SD8Qf/cKX?(0
fe\L5ZS8)=ND:;)(J(J(:YWHa\FV.46]704SQAM6bKEH\C=&gD(WQMf-FPfFKPE1
<]J40W#^:29VJ7;]/<4SNR;Z2-LKgaP,XQ-FJ#;@9aY.<?@/,?7&6899d2]Za2W5
F,4\/O2774LYa;#6I&78VRG@C4Pe)>4+-cOV#<Ng#dgC+P6_0d@4)1aAL\;We&]Z
dfC477&[;8[IYL+KC@<@7P#_4e:e94)P3;>5\V,D^<O/9X_P\X=Fg54<a&\fa&T)
C<K@SSS^)0g.=L[V)JF&N87\,&Ob87dUfX5+Kd?#W:=Q,KA>\WHJd3B3gJ>)?FWV
F29d4/IWNT:4>g4a<(0C(=\VEB.C,CY[>#9ISCf<B3WS@T9=FA>;.69ULW[0:??:
dLeR)QZ&>\<[Y30G6Y,+N_8-M01O#;6Ha_M#Eg2:2<#-BIM:>5M:aW5,P]bcV+dO
W:]dI=U\dUgf(?gH02D[_^T7=GRR@P0bUXa=GC-W&JM1VQX(:aSfXc</UC=\6C+?
#,d[eQ.I830a.-0:-ZC&5F:C>P>6?AVPNggd-Z,OOCL]BS_@0R</)4U0PDYab(_g
48[0=\B@Q1N[Eg-I;ceFT;<8MDccZZ)cFg;-QF+YVV(S5UP\e?BbLbB_W;Jd(63>
>0LMVSVEIO\V&DDL#7-NQF:.,U[@,F.BV\Q+J@]540FU^EeV_@>=Gf:6UH>G0ZXS
QBA)&gMFVMACE/?)cY8A.O.W[T.g0@e@5>IWR(#M@f)/MFORAdG>4O.[-=2#+51G
_7O>M+7C8IV#,<SX&;\6:f+]aT1Ce/SJGe;1,I4#KVU.IOZKgYV]GBdf4(R8;)YQ
EAaf<XUF)0a7C>13Z;dV9+H,?N<T#5O.7I]&d&OXJ;B,<1\M1IN0J@UPXPQIKR1Q
P@fIS&#QR?9]6.4>^3K]BALcPcGMc8_b]G[:BFIYF?GPFU0P_A&,\]NQQOG<&FZA
,,-EVG[Me4Q[@2BJ]f_L9M[e_J<5FLZ53N;WUXD7ZCDJ&XUQOZ0@#/?e#]97BA@J
dL)JgSaefABb<BAdf(YggI[E+RNFcYC/bYO,aDe6We[2X.A1R(8&>+/55B5@GFJ#
P1=.YM\d@U^R7O=)c?A.<6Q2[3^Ab=7;5^5A;@.ZV6U[_M7-(3E5&KE0O#>A/(^e
>QgU,_=QGRe(cG:;b,N.I[^)H08eH])U6-Da3JV=97@?Q^-76a[M2I5HOJPW/S>Z
fWOUc2T@H4.Sb/PV<VJACBL=12\:X?:;A2,ULHWTT.c^TU]YS+H,96P\YK-YJ<1e
3g)+8JgeN&b:O36O&#^:S>K6M7eHM,;b,A;U]?g@FPAM6_C_6J7cedUH41:3M2+R
;#1ME2OB\7Q/;(5e8O#S.b?XgCYCLGX05.J_TWW=[)[W@DcWO:g.].D?JW&d]2I_
PUc-8dQeBc&eLW)[F[LWTU?P7:-908A>FHNB/&QQWgC\2;X;ZC_=ET=(O>F8RD,4
H5H/gL6\[A=-\C]^G.1D;7?E-V5HI54EFF702L>f/Qe&ZOa@cOHd-J=F;FI)-;TQ
:_3)/X(U:TNBa@&_C#e(;KY\ZF\78VNP</43aMVAXM,ZN:S3RCb7?FK:&<+f4N=H
bYJa-NBBJdS.bLX>0(JUcMa?=]fJadTI:0bd6Tf[\QJFgA@3_a_,;CbGdd9gDNWW
ZA95@S@T2K<C=QAB8Z;V4<R[9N4HJ2AB\][0A-:R_75(2[(-F[L3/#Y[(]1321Q?
YPZ\Q)f;R-MJ>W<Z+P3Q[\]dg8))K3@B<N)CU6;?U&IZ]JX07#CW(1I6bXcJ#(G0
<1+&)f?c9]);,=1?Og_03SM).1[COMTD9<+D=Ff+4ZgDPfCb]@Z.P=CWPY9WbNe@
I</1bIU)[0^Rfc5\W51N)+R<YcZG:^F21AQa:\?KdbF>:_I;I7Sf6J.Q\F&H=9V:
1--^K1c?1S[B2X^-_,)M_],eP(6/V?03][fGd9=H?/L27TD0gWf48g7.]Of>>6T<
]BWRJg[\^:E:VFKX?J/beJXF,MH5edcS1[4\I4#@XB(P#(g0#e^7dABN?:bQ^Z.+
eR]4#Ce;DFd#gdUM7B19II[d@&fM2,9F)Z9\55E(N?:@L#Hf3K1(Sa:9]GLcP.;g
Y#W(\P4&>ZTeH@K39eH(1/eJ@f5OP(Kf#-X/CR&??fT=NG<S1Y0BFTRaPR4Y0cW=
dba>E2]K&T-MH/?D975b^V>c_;=K&+)A,6@6aKEXgfeZP[\CYfG?a90(ZWd]=X(@
A^VS+Z83#73K05N<.5eP\&Q0@FSeWXe5M=Q,P=f@155V3VED)E3IKcLKH.P_OHB)
Y4KX-[E:M0^=#ON#&4\LI&?Q/.S#&PP644Rdc;A#4NdT<QGWX23f-FL\-(M_;4@3
R/JSOZWU^bB>&UbaE#8Le^WeI-FGD;-Z4NR/9N4_Z+O\S7Eca:3H_P@4@YNF/JGH
e-E(CPdL)&4P/JC7db&WXaHL89WPK\&#J?JdG#@23[^PF2?.9K\-),+RNZTJeF;M
E3d]:Z&RBJQ.VL&IE8\baW+e0=:TCVPKIF@U@BIa3&+X1Ab7b&K_,,P]][=0]\9f
RM48g>BU>1DKR@]->@d;9Wc;faS1d,c5b_A1/BJc=/S=60&T:2f_>,CE-YF#U7e\
\/2T>D(4A6[RaIb8dBEb7J&SQ^<^e9WLg2&D,5S9Ea)/EJ>P:H#TBCdga3f13JVg
&&Lgb+DHA#WAG<#H.Y&3d_S]-4V7W6-(6gO^c1-ZG+\#9c;8d\ZeP1aVF#AP[\^B
L1GPe=6dd##ICgc1B]S\M\,/B,a?AOT8<VI;g,f.?))C^JK2Y&f^4)e6P\>QIYUf
(Xd<76@^dJ)U62dVSA/df;&R1Pea]-gQ2XbTG^\)<)^6H24D6,&CW[d_HZ713M[N
C-\PBYN]5M8:92+D4IRIc;7&14IT;D508J^/2gd0>a]Q6+d#?05?9U7YUdM?,+PK
-gf;\Qb]6+M<R#;[?S8e0YdZ@SCML/E&TMUH=.0.[G(D/3Ca)c/.@<94GM_eC70:
H54B9/\->/#H#?a_WF5_:@cX+31UOJ/C7AN;^/2VR2=I.;b.eKIC=QYH(QQ4@JJ4
G6Se3B:K1P50<IFW\G=(Sc#&Pg:H@54E6[cK_d)-MWW^^D7F>2U3L(R&eWN#2We&
gA+7\2(F-)&c\XgBf&TE]]UMO51T<E,;FT;#S2IL>2:YGD]XC4-aST&E.9GGVM8M
;:>d=XQ<I?GJ\O-[HQW4#(98^[JF?H_IKF>=W1[E+?6L),KW<:34H5;U54\=<)3[
O\8Z1(,ZM2@@4JX8-NGZbJ1\,BM/fX5)=7_J<\)+,5@\/\9X3S2.[]2b,OK1HF(7
LdMT/FKg&RV6c?]EXTBJ+f\BIHFYEJ=\-K#?G^3[X.:aOZ>U1K6ILV,;/eS8GB3:
@0U?FV7dBE,?Wa-RfS/95+K#TH[>10OAD(0C845?E?7a]_R7T5Hea_JLB#AZN_=A
BN3eZE+HQK&dX?13C=;F7JPEfW[2fO.X]?>0\f#B-?RF@<^\#JL=+#:Y2&FEd_4b
/3-CY]HN#a&:C2M2)#QBOfEWZWa(Ddf1C)2bOS8Q6TZ3.JW[V..6CVUP^Z@J1cHA
0/aecQbXB1T455W5^+-abg&:RY7ZDQ#R7ZW?bf(6Z,5DZc#YL.,HT19-4N=U_g?9
RDa&B:S7Y\(V3BOcU6)LWGcc??&Y+dZ3Qg-ZM6(d#9(--(]WV^.G5Y43I<cYUYG@
Y1U(1]^;68U;Vg6A9Z\BgA0+N:Kf/YLc8J/bPDC#a#+Yb?3Zf&E0=e@cMT9Q^V9C
Y/_9&DKb072YZ^&J_V/T>^:OUNLI3Y/-R]T4&BFc1J:VA18A#^:3GAeA&HT5_/ID
8+#?_5K-MaQD<\/W<[(DP)Hd@/7?KBUW,Z3<FdAMVY5M]e=Y6dI4GKb;Ec@U^Y?Z
O;7R,8-Hc@D/PKS[8DY=0[SRAF9;M3,:@0&C>-cNS(=<Zb?;a?EU<(P:)e?-F3]W
Z.;G1IS?BP2LePCNSNM8I^gMP&6F=aN@R9EA2SEDV^c)f,0]@0\@F\_g,MZ8/-P<
LJJH9Q,BW&/XXS-&O/6#BU6LL?Q.eJ]9_<ZKeOb+/CYcK,(>Gg1;179X2C,3)4&=
VV(+C?)cAcF6DYRZe0KGRba+<_e/U0(/2MbX<S=53F4+)XHY(5Q+J5Dg#0[O=8T\
RO?)PEUAI@\CA8X2bg?fBTVR)G9_J7@WFRfEZ<<CUdB@BC;\BK-MDSL:aSSGeY+<
9?V9F3?#70SKWQ\H9MVNADc\.=>LdU0>\a]JL?[?_H(.C)GJM[1V&d/E,eBVcKC8
)M#1]->g?RN74_Ac=dcP>BQ:bgfSL)B5C(=4+:Rg?e,S22gbH9RQ.E?:R-IDgeFe
GgWY3,?KW@RM?B#-)XdW+4W,5:K.9^6W^K)@(4[7fINf=IbH_IH2b]YL6[R&]F]I
fYM,)<=\8^1\_Y/.#&2IHS-;e1SDH.#L9C(SM#=)/Q)U^MPI1(FA]1?7-6&RC^LA
g7WR8B\\8MH(]bEP,5#:-CXa>>V\5+VMaXbP1e0:#\[-)g5COG\:(ZPe4O?<eC5e
/AXJK&OI\R]90>Y\M&8F0[(-_Ug)Y\V-QB+\.5/dBUPFQg,(@BNcWCOdKH^D)C=+
5AW/>efHO0HXe\bZB&<eUeDG2g+0bUY\SH4/bCZ^Y^2;)B#=.3CIH.7:2DR,LTHD
EF8LFGH>R4RQgK5U@9:XA;LG]JS>+D.F:G-GcNOB1OfXJKNK^34JTZLL5eY-/W_E
2DM9V]H2K)P5XRS?FSeTC3[[5(=)=:OPc[O?b:N5]ZI>24(2QY2f\>>T+QD4QLUY
dFQYRT,V63[WaFQ1A20@UBT#>_cbJVe8K7)a87I5KYb.e37>SD1=cWb#TcEL<F-3
@V/+F9a:c57eWXQ@2&L,&<88]Hf=U\bOML0#I@;W2N:.2H74ef^]:/#+IYLN09cf
WYQI\b_:D+V>PATY\;HOKG-\&F1,S)R428))5]:O(HWCA.RV_cCUAI<OO)YbCEMG
&GC/E)&6Y7IQaaV:.g;,T:UWD(X6/JQ2c?EF3XbBSBI^25R2?.1V)dX[R.R53-)K
.,dYH[^I/P3+\cb8+(CA=]@Y0AI^(R-24#6F<CaY.NO8+e]#Y9a\@)Rb3(fKFL>7
I5X+Y&P(E&CB=H2;1R18&@.CVUQ7d@EX)dO;^90D>]gZ&1cJV0e,ZDY@]5[P:/55
E&OcS-SREb;6VH04LS,#<;gXUX9R/Ae#aWD^#SXTF4Y@F-a2gQ<McaS)/aVK[H#G
261Y;.#7:7:)<80]c-T]EMN7_LZ10a1<<>ZaXUabV&fRJP-J7e9(I^)N.QeQ)Bad
NHSO\6WJ.#X;VC8T,/5HFCbTK;c3^W^:V=Rd:2GdQ4a+ARZ7:;H?WJ5XX(g0-JbU
PGK)]CRa&NGQX_D8MCgg4:8G\4JbX::8QA<=^5^:]b\E9)YY8g^,KeHOX^,Va#a]
.A.QbEC_fbK/2]^.c8S=&3),KbW@+[Jf1KU-KIG3(82#GO2L8#VD5[fNCW9^a4]J
?Y^7;0Pe,D;C><))O5VNFFJ<^NZ@[/UV:eV<>gB=@-Ng7.SZ8_a;.T&1KF8:IC52
CbXJLcR&@;-[9?Z@#P#QG6IZ(0>QZ+4aV23g:aa.8F3?f@ADA[:N4,I/5ZEfcJ>+
\YF]0g=3YS_V;^:c+=G??Z(PG\PL]QU@gHW=(]T.T&^-#]V1I,41Qd<VZAYOKeDD
b5IQOJR5JeM)O-SI?dg7F+Z+Z0^DH;W+4:[VBWeV=U\;a,OKe)@cHdREG1^SG3S6
)/YMI]7ZRUM<6Qa&@(/Rd,#,CMI[Q;:c2@^<gYeNMUg&;L[NS#QL[_;ALB+VgRDA
8b&5(CE?Df/)]d;aERL-JZFLeRIB[2g(]Z(C\D-Q2W)9/f^ccV42P7K]NDD)C/d-
NKB,(GDY#D/O(-Yb5FO&,&:)U<8Z30JJN.7JG61NH+ZAPeXeca:5H#BD.WI>FUe0
--CEVP+GNH@2EJQ/e>+4&X9GHO7E0E#3Sa94HLX[_1++/#OU2U;[&ATD8.B9Z?&E
MSBE7[5OLdCF;BW58VCJAKXf[Z9UgY4WfT_K8[g_0\B+D-0NR:dg[MQDb7#gDcW5
R#W>P+0]8C+A.b^P5,KJ?8IG5FW#GPEaQF_-(5WVgE1]/H=]8dEEa+U\B>]JgYX(
^^HF?<0QU/SQ\SKXR7.E1.GPf0;.>L_MQYZ\RQYJ9aT/X5Mg3;5-4]Zd4e-XdD.I
H+HT,Q4b==eCY59B,_IHcBf]K#UK_J2?/G^-Q-+.PBb9O_M\_(#7QP_P;U^6/.B0
(D+Td7W#1SE#]5\5^&]&W95/b6g9&U=;\d<4,/8d1UO:9JYP0U/.LQV;gOL>a=R1
])G^:<&[CCQ<Y.aV]QLE51X3.D>6BLH>)c.g5(d1bYbCL4Q:XKT9OVTZ9bXZ4?,F
3H&K(7Q22dcKY_99bH(X/B;T;#6Vb+_=O5+XX?RDId782HWJ48MJ47;ccIa1@1ZA
ZO]7N@Z0<LMBVIa0:8c=428J[Tg#4/A/0=)YQDV1P.L<V;_)XLHdG..S6J)C5DbV
]+THVJ.SS&/])ba7S\2SB0QM#)#Q1;@4EXY4C#_F[R.dD_6E:XddL<<MP^\2M_N=
^1[A+YSOUTJ8LagCPTS\c7Tb-6NKd^F#R?-R=a3]U_eG)gV,6(efgR]ED5U9(DK8
?N8#;B,=:Y#IVb@DHL-CbW.K]@f>QgQ[/F1:MbaL&_^D<_.EVCeKYN<e7aaZ:V4b
:KL)TUL2(_HH[A:LQ]#SY3MOAgU.O24\a4N>(aJKUOa6A/527eNY)-[@K8?:G^c0
X6JO4BY?8^)MCGgIdBW(W#UKC=&]dgaUZOPgW7^F[H5c<b#A;+3.-W,JL71LMb47
V@)&T9&S-K09f\AV\N_F/4;Y29)3O]d],0]KX)4b>_Aceb_\.0cLR^E<DDfDS.+-
L,,B@06ZYB[H0F0U)=?DZ=WV91_+(d2c&&RgG;d848b]:A^ZL(Q+SO?:Kc<-;J&>
\TUM1\LZO#0D1\9bG8==feG<d>5K3U.6:aWV]P=0TKbIC2;PTCQH//LS9O\eCW^I
(QXGcG#g?eFKa24^=.c8/3OESD2K@Ad=JUYVJ0:9]C6dcFG6A5>VR3-)_AMFL.3<
7ZQa+S-b?>;3X;U(-]E-TGbD@V\gR8^PG3WL(g(]4ID.@7aLObJAC[?0VR+P4&6-
Y-.:ON8SEQQJR(>QYfV&g^e@2c>XI,b[P_X-YCW=Dd.]?A34b33Y/UCa9fXdDU1J
20=.c7fe>&3)+#A@(EdSJBUL^8F3_187SSAA<S_353CZHAB]RV>YTA/TOd,=(Sb[
GQ>(KE;6B-=58>J:27Y^c1^/#^SWU/=69Rge)dZF^7^O;dZU.ZFO0eWH((G:?36W
W:@Dg]/#N<P2+O-8(PG18432M)c:<XPYeXJ3#/\ASX8d_M+8@T9KN4R7_6_T^#aY
>MFC4KBF^XDE&a7gSK.)LEeRP[^,g,HSD12CV(B>cXJ6bWZ=AFdUIB8E8S.VB26a
RR+.3_,?U2YZ#^V&@g?c:g^f9;a8?\V+)#9.8HSPc6U#7:&+Q(2@KWE.#+R5_]Gg
QBX78SY^b8XD46cHL4-9JBe@=72gL?FEIJVPQH#:AMP.F,d.=D8QLG?.Y;C5^g9-
,0\IG-4g5.-3SQ=,fCFRE,&6L8O2J-0J:)0B18dWC0))gf;d(F^GY;4?7HgQKACW
6e90:;8L9_GZK0-7SQbR8?8:1Y\P#+.Wg;K2?>CRBI:<=JPYI__4;b>RRX@f-HVe
PL1Q=:U].(XN#AH/3#_>8XT6E3RR.DN+eKH3Y>c(SP.M[;SP7^97]67T:=TN)ZgF
#d85VYB(J?DK2YS@\MS1#(:WXaU&P1eI&\[/6-Wc,/S.O-CE4cXd8[a0)2[2>I2\
MBC,J4GeN7gP><c4VYe/>3<=&)JF?d>+aSP6HP,7UDF1;:-AN<:AU3?S&-.?7bUV
Je7=a&>#1+]CKF\T>[f,WP\_>:M-/2b;^=)e,/fUNKZXO&A:LgV&DDJbCeEc]^=X
1d7P7IRMHETd4MV/Y_2TLW<O7;<[,VW;Y3J3VNTW^MU)?OW3e+S]3O>GHC.2EW_6
<>4J7&IFS@+5DF8R.[Q.G(FO23cP5g,AWdH_F^8JGT;1=U]OTBT:O)7Sb\1bZF#2
gFBeZF#Y@g#ER\fR/6W,O^QY3)MHC0P;6S8fb&N\+E#:WX,--57S>&-H)>\b2<AV
81+7DdM-ad[ZBI:OGS0&K25.P19&-f)_OEZ=KE#<G<)1TZ3F=(5K0[VC0(^b[Ge\
[\\N\#4UKG?]CXZgYVTD0GJAV\>d.@/d5_@XF].#Fd8b@g)O20T28&LR_O(\[IU9
43:58g=2AAIKJC];Y;e2FP0[3<0Vc(;(B;Q0;XVVQ2B;9c:\WWE)=.NC<6:@A]+9
AEQNe?DN@Q]F7FE0c\G[FCV2CH<(=G]1#R8-&?_^UNX2+U09b6+&U]AX7g_6=\0W
4@.e,K+S;_FXWe=_)?]X,dbg:&B8PR<//5TAH,(U/K9J+6F^VC2b9bIe1X7A8^b.
YK_]ZI1_SIN;g(?\_.^ID(H@9cL<;]f9UB2X4-78HW^NB88)>@aPObY]=0#fgg7]
f/9\ZVO@dfH>]JR+_0HDTUKVW7>9RBN<La8V?BR=e(+IH.FZOQL#<J-<OI](eg;,
fdH1>69OF8X(Z(1a=_4]ER,P74+-M0SS&,]G5eYR(G14/_MGMK+:TeJ)&H<E_#Ge
G2O#.5K5VcTXRSHdDKT:&VJFA1/@P-R=2#=^4NT<[0I1e_\[bd.3eOMEb(=&.7d=
6a@3P3g0K@X7B55SYTc0H1)LRBfAE87S.cI_[/gB/KZBd+TgE\d+a=_28/I&#(P#
75?EK-b]JdMH<Y,@JA=F@NAHF^eIOG9^>RJCR-92@L6>J-.A,3A9(d)d^J:eL/SB
DCHY98.RL1>.SY@I)9BQ>NZWg:@D#,9bULI?d=45E?W?OST<6>>HZc;^0MaPTRTf
.YA-af#fbQ[89O#,FT:X^9Qfe6QH2K>;aD=>6#L74Pb;V)cA_3XG[S;?JW;]8ZbA
&GU0<@<V\YH-)1C=OaaJ3OP[9d;VDWa?W)Sc8](HOX+GD&+;S<f;J6>@CLS<>d0E
5JZ3\-JHA6]E\^HL7_GKQQS-15b(W\_.0>ICX>BWAe^7+.e-[:=_R^[[K8<S4aW/
e,Z)P[PMfgU>,KL;&L3F0g8fFQbgZ.4>E20g9G#P0FZ31b)d,U_(O:IR=WR[>X+W
@dAgDEN?YP,b]N,[4[\B/0g4e<K_<MgO<)^VA3BEMZ&Q_=WJ@f+1GYPC?,EBbKaZ
a\Pd;Y:I==UKXEEV;V6ND^B@TF257KZTZR,b3gP,X#SRA,C:f\#cI+?TA&fNg8Z+
6S-ZN;^8V5@;f;.A0cBb:O+V:^ScV&=:d@<X&B=/gCTY@TG,.[b:?JMQG>0;(b+Z
I#>g,^&GP:<16#@7V7B-c4.;cX^A3RXI/9Fg)eH#ZM4:^.geEK\f(=,->-6gK.5L
:V+gQO<N:NbZ,eI2/_\]46=1K3e_CR(L7cY6XbP\3<LU>>I8DY]U9BK]_La?WMdR
Q[NF1-LI1@MUY&;^PAL-QabfgNcM^I^g]eM4H?^ILYJ45TDEPZ[\d>:TP<He#cKS
cV;C.Bf+3E9T\:Sc<,CR-AefVFG79KMdFXK:<.YGPf,c+R[BM2[58MQB]_[?>-L1
QDL\]>fR>Lg]8-UYQ]3E@H;(B(b(OL3C)ODF]]AKU@-WGgZ<8Qg/3L.LNOa4CZ_1
L]3)bE(7A4]1QSe_U4a4L9;<AcJUMg1S-X)>I,P:W5:D>f1V8TeKF,Fa.5-Q,.0E
DLX+WAVgc/\1e411EWH.OB-0,(;];PT.L:FW-\[dfUM@(;\#M/UP5<^4LZC:SBUb
[RDBVd7Sb5G\E903?BO]=_cd@UF82K9^_P9/F#.fRd/[7^/J=IHI#L88B[/LY<aF
:[L)2[FQdQbdK=RG39Q&HaWb?3C;,V7JCbUQQeT.,c:PLK_=7;9H\7Oae+S;AW?N
D147HOA95ELL<+d(degMf?fIb5Na9<-S?,ZN=RTeY5ZOT&&RFMCD#.\D4?J,<L3=
::N,DT;BR35/E]GH)M^9VMS\#H_f/LB&FKG@\AV>Sb>I@1Q6TKb_K+5RY+L;V1De
N&Q>.RgE-HI]P^+)H8>^WHM:D)/TDDH(<#)F&dIVeTd:gXT)\de[aVVX1YHV,A_5
&4:1^bg45NA&g6\NSe7<aHFg]ZK-E#D?G+,:5Y3]f3gB&dU5cW2<CeGUaELeN@P,
9VD[MA=RU\UCOQ\f]?4BWKV:4OD^)R#OEN74.4ZEA+LA;KB<5XQ<=1MH.TJe5bY&
V5TX0-9L_[3DO,EfASIS1<QH^B,D>+J;<\_H/)XQ@.X8f.Rf^.dWR?ZL8#\@DX<E
_aU@8#eXB])B[X\0^PFf_#(I<3,KB@GA<-Z>5O6IV)\^d6OB\g03?H6\XW[<K>TY
3YBKP#KNg>DX2G(1;+8g5CO(.M4B&10NeF-@CZ2@HWdR96gZ]1PR4LXTHKc6O^KJ
:Y,#5=8UFdc8G_:O=650<)Nb0C?_b\\ZPE)TXA5-N#;PR#Z\&J/;dfH@KH9&Oac]
..f^?;TTI&063WRF1MbJU:TG(_16=#1?+1(I?9)J9dG^J[Xb&-^Z#PcH1e1CfC-#
G]RVQ.CWb:C4PP5d8LBW^&PLfE]WE,RMNB)GTQY+V7Y\&3-.B;Y_0JVW7f>Y[g+5
GM8R(WU1Ia4#fd=S?;1^8LK;(7&gXWK9B>c&]^BGU2@K1NY^SP^@1JK:EBeaD\d=
T.:#M&H34W]A>U,XC+5F^=-d?8-LD=(KfJ/?=?98^LY9ac5X2\#a<P1[;C=#Cd7Z
+(6OM:-GE:ZI+\HS<F&.bAe:X5VSfQ(:La[0Q37Q=bYH)-+Z3KI5=,1_IK0##P#4
&Mc/d,fDeRO+RDVZ+,Qd)DKFV[9)P0(-AW=(7_VWM+:^WBZA&?D))2c:9<5+#dPO
RF8,H\ZTL0WFTb]cTc:))Y+C2D48Y)8V[YcB]FIfYaf][DGQ(K>,_e7EHYI\]4XR
E&V+:.YfRKD0R[J69_e:<JE;2/MZ@G/+5)<EO\,Z:22IVaAbD^2#08a[W6D^7)/;
71T,4+AI1\2d,W;Be,a-&_J8Q7][DB8^<Ge[^;\P<CBOKePG3/eAD5Bcc+NO[;;6
8HTGM/J4^d?BPc+_Je.URHTK?c)cWYUE++(E=fX=3;C<4gSVCA&FV4)D(F<==U16
cTX]^OL9,bWLNK.-=\BWTf[fIAEP.gMe28YAO/KSWX7fZ@ecR9XZRc/FVZ-B77Ld
ZVL.6(G/<]ZYLJK\X:2e4UV4.;W6-_Re=9g7WGg;,0ZJFg/\GdRPCdb;)B+FePb,
@JCO^C]E0=N7UeA&M+]Ud8?;FEeFaCK]_V2JdIZ4<FM_G70YY2N<9S^@#/NP[GB)
16DY0C4cPJCJ84#cBHa[/J0a&R)1Y9Vb#\F+<?VQ@-_YKY>:;-:B6#?e:ccRe^S?
@MMX?H;GCf2GAb(WO_)[RVI)GI.75=+0e9_L,2^SI3N&dRH9<&?O&:@:N@bZY2d(
6=Q-6Q[/LFTS]FZ7Sd8ZGgI];cSN@Z?]0(SYdbIcOIW)&DUS[1F5W:a;3<TV4;]K
ASH0?\:F45.f)(]_X2S.</(5(/AE7G0I]f[\/d^)Pd0,77NJN2+A\e3P<?dW9L6d
;OY,&PN_LJK1fSDC4#F6:IA?;R<^^g.0Ib1)a:^d=]&aaMbICeU8QJVL__MC6V(c
8IK1VC#dM6aX1YGeU0QA1d](aWI.I9VPa#MB4\N\Gf)M70QG6D8#)BbUIg43Xe38
;LU>;#=#[eKP+7a?#4bAC3gS7O<5f]&^4Jc]b_;UI);0;C46G9W4=8L,82J9)-Hg
S@J,?O[NSDFSf=N>:AJ#6dd5g6U7HW/)4/JaVf#bB6;f0W>56L75VGT^<M_9V1Rg
6^/\+KF6797DK^QI1XNDba/ZKAMCE;?:>#RZe^;eMX@/LF=E:P4U431DF//O4C#N
CB.?XA,bTSc@#55L?4dF786/]F3U^>)FCf0N5XWQ(L(C]GYYGFA8A15S?3Q^>F25
GDQ3+[e^M2:2X#<BIa]<SN<d0O:Y#[e_Ve;C>a/)Y,RfH/J&PZ>F?G&M.cR3O.Q&
OSM:cMaDY@dT8BX&212_>bUX#+9TMO?]TC)HA[K2-J,b9#3HC,aJKN(78&_bT62[
Cc&c@cZC#O-@9-TJaZ[D<;(1KKgNV?10EeAPN0K(-P<+5=NPE5+]1c.4=D\GP\8E
42)D[5>@6F(5V^H,+@RI+J.CE_ME92#Q]RRTaVA9IZb(eS&XE;EOX(>1K5F2U[OY
@Kd3fS.=4XP18Y;UeBdVd1a(WN2,e<3#/bHE,P4a(+:8Feg>cGQ9e?aJET)V4&^Z
?:Ub\QQQK5QSA1_0GF8C^.H\O+/L72c5JI#KO]5\G.8B,=HZQXG/;1J=A:I=J0G^
<G:J.W1+VU1GfeAd/O2,]K_/.>d6,cHV#ecK<+N>H0^V6]b#6]:GFPIUYP;Kdf#A
MN8SVIL,RM,1aLPZ=Z;9F)+EG-Ag3>A\\R=9TR]GCZ]1b9;#XWS;.,_]8G#c&OTg
2A6?D:293(<WXB(38=b,Te]MGd-2/=)TcCZA@CY\Jc<US]g&,=&eLd4FfW&9EFg.
b;#aU3a#E/Q=B@>N&fLIb:O_<=0<;:0/^\WdcL8F#JNFdKa50c]RGg0C<J\E/]L[
8^>/IC\\C[e&#)J_1G;A.[H6HU10,.FG@1#E@&/8=K^Ic&gXW4/Q-5M=K,W[UK2S
:#dZO:a>FYCS#\3XH4+8b:=DR@gb2?4LNOQ//Z2Wcg\@fZ?(B4Jg7/dQU,)5:<1Y
9T/K0P)#?9ba:bOIFPZ)<Bc]-]?JcX;D_U(\B)AbSE^7P=23JUBCMIYT6O-R2\e>
7dES<Q(@YN)TDP;10@8ITOHWX2YNN2]E)5dY+27.]_Y2))_eTFM(92M?WIG0-BT5
\1XUD?P+e5F-7+)G??YL:JF=a6AEa]M:DVgaJUO@cK+2KPA@Y:39T,eS)#A_>K4[
f9TM,LQ6-VVFU0QNG6^3PcAHf9+[6+gNQ7JgRY^)3;@aLA:ca>2b,@#Q6<b&4([D
ZI@Nf8=^MS42Lb4cN34&dHN045X039f8+)83ZW(MX^fVRg,G0Ug9Ba9>#SN/.cVX
6V\U6M#_E8)8DGI#[+-RG@G&??2L]T\WZ[S,1=J8gcC:]/0S&_WA-GK>O)^8@Y7@
^M;T6#gTcb1/:GRZ[)6HOZLU^2T\f_#WF0SEF?E,WJ.[M>3bZ8)GJW#?C\?M_Y:M
(\)DP2c9Z39M[c6P>1NVW4+;fL@J-UMPT/3+b(81c/QI?6I&,B8[M,1_#.F^E,Ma
F25P+\#Y4768OV:ULD,TbG;e3H-IA(WM#VR2]f;]8,16?[?,d:(/5FIgB?9WdVDY
]Q&I;0S11bC:(,T8+=)U\HE<_<EZ]6:H5+CI67)aV,Nd&NK9CWZ3XBLIVO2;.gbf
Ia6@T,(+.789^:f6P.2VXd2X]&J];]=V(KFVU,ZS/W,d:]U9UFAdIBIFEC,63Rg(
Qg]H0:MgbSBJ]7UZfa,SFF2Cc,R3]eGWb7.d;3P@/08FKG:9&SIL_Ed:S0]:_.X.
;eWCeZAYHQR#MWa\1YZF<>,YM&LAA0.[,,<5PR+54Ef8=ee:L.C.GKLZ->\?LVQJ
OI-&U[(0c609@4DMBM;LH]^<gJX04#&_D/GHTV5R:Ma[\T0=-&_M((AVXN.:C[:6
HcR[U7&XSeeIe=(CQJgK]W:g[;[DIF:BNJ<#+T88\[DM+-J\N\J@dZMTPQUZH?)/
C7<:Q5=F<D70O(a-:CS0>g-GC?G+0F2)P9&)DU#)K16A:9T;>D0VFb-2V9[=X@+4
-TD^9<.PE2,Z(P&c7\WTeXU@4BEV:-4XD?7aP=WL.F6bM2=I]31=DDYR?a06IL0B
7Jg[R;19e4GLTQca=I6VBS.5G-&-C5-MWII,<\@(AIB12F<VWR5ZE)I=;O43YfGP
TD_AfGZFJ(@EcfB^]@\Y2bTPWbbG@>C6M\;.?a)L3(L\G+gf7K-<]/Y4N^+V\(4J
]RJR?A@<_dcI&:L4e)N[].TR>c][6]S+/_B#97SdF.Ha.0)/2HIK:^0G?YcICRHO
.DeD]E+:CD3^WMc#L&6Q,\[8_L])C1@LHf24&VZdPOF?LIIL(7]R?]QX1Oa=(5-R
M.(S7W&@UEJe3e.T?M=UbN1K<T_3cG^17A5R-4193OS&T:PdQWID]K1Z=39Bc/?O
/R([JXCH@0AO9)K(/f.)bYD50)7JfU00VD#5^c-[;]#\^D_/=L/<(PJCCC=L/LNR
]4@N^d8OB<0aJSeRN=K1dW)(K^dcNJ+;e&:)MXV2,ODF=Ea6:cECDDa0+9\G?3CI
.=U^O5ed@XfHE?&Z?FL[Z(]6R\aB#+RT8#JMKFPU]@+=RL3UWI&-UJ:IJB51cd)8
UU80O3e9AOc>OT2fP3F[?_::cHOagDG1:2J:Xb7dS35c>38[aIG>8(0/IgCbc<X0
[BIIg?A7ZU,JSJ05<7b().]G]@@(4QH8ZIeM++72(3V+b0JI7aYN\DBYe4P<.:cT
KO)Z-9@XggPQ]\0JSD[O9_6=9:)LQB0J)0L\VS[fB1R-cU>,8NDD=CLUQ.]=7KT2
&XF+A91HY9)BNJM=22YA]S=^8P<Y6VL_:H5WPOOfWTS;Q&[FD^5KI<#CFM-NG^HI
&U],eS+#CQBHb62,.2&A+_DeORJL,S;eWbU7:bO;&TUYLAG+F;LTZN7&^-H2c7&Q
0#Be.,03ML-N^:e:OSTU;S/dZD,g^GL\=dbR\NPbYO+-W2.c<(0TX]+0Q=.S:,Z?
4FJNZ6+@FMNaOcP72Ad3+(5QTN&#-dQOM)DM:DV6:)b\I+8Q&8LPf2,MK?Q77RT0
-9U:U..MF>MO,(=gNcM^.;[#^/eM3N2^=T>/1=_FdANN),&@X5B\,:=9[T.6.=Z)
C]NQ:&4gWgDL[(FdM@9Mcg(5F?\-ec4ET=2N-V<,R.</Q3a5S)X&POfQg?+=?<&8
Ob-:81DdFG1W-A=^H8J^:O5Gc@:?[1?aQS/DFWXLCDd&J[6.fd0]PX#HBS11MCa\
5?KQJ^ON,XEW\F.c[H[QWbNcAea:1_71M2LYa@Fg>5a@@a2QL7BJ_cGALB>FMd1R
F_.]C<K9M-GSP<O3.,G-@=,gc3Ef\gG7eCcV03S>\^5H+SUXc<F>F#&\J>3HQa<(
^61B9SV/MI8HKRO&ET:MP9eAbD>U>BCUO+D1W>5+BTDF;WO=9bB0eNO]1NY\=M47
RSM+VLLZ-B3gfM8Z17AX(bR\PT1(>O<CCT/LCD.&/8P.2>?6b<4-VYQTL,0eK67Q
M,R#)fOX>BRCQbP2]NH^4/C;V<^8157^&5c@Z5Z-]6ec-G@EJ_LIL>;gC[\5PY/V
TbV2+V^ZWJ^)5-W]X7K^.aB2&FEQ3.b/bg-cddH1c5F2O-DaRQ#[FcgdW27E>9He
WEM5[-UVMKb[^<e4a84=SW3U,>A>4=a)a7;T@0Z5dcI7SW?J8W.eb7<>Q3\Z2ZP0
\IA>6a/_^W)B5DeD1WQNGQGBAE1CODCQ=6g/HBV[93V[1c0c#]HZ<@[RSFDfQ?^=
A#C7&;gX_#9[7MIIe:DEcW+4B-><>&V^a/#=;F-M\I)J4&ag(U\CJ,3(?=)K&TOS
QY^R/RN^=Q)LVJW:QR;1f5@LT1-HHb;3GCHad];4,OGTg/5;/&[aX0FDO^_#+SQg
;cDgT=EEc+(3XH#Mb>4:S>1R9c/?1MS5R99-MDAMH;&_[].TBZ)c20)#]XNbCaL_
,WNVa29RS[E[@D+49T/]W7KTcTN6cVePC3Rc+:JD]DT:3;N-P2?Rbc6]f)bI\?&#
#++DW6=A5@F-;WZQ>:S07>>?<]87bM_LeY)gW44=WN+GC#F71GMZ3HddAHV_[S&9
/0/_ON8OC/^S/f0+Mab/:g4V<dd)/A(Sd>:1)a&??.X3H9\7DW#W@UK9b@PS-[?9
X&@DDg:=[P33\BC;NGaH6?5/#LVWQPZV>A.RSf1a2g1WX?C)[25=E2dE)D;c6D(@
#]^EUTCKIQH>[&e0=bRd#_,bKT6U8F7c5.CL#@SSYJd[8PJaNUf[fY0OE.7bBJQ]
M]&=7A08]1C]/^UC8?@C&2E4e5I8+/8:W:7^+ZNEQ8eRZg>B?^=g/_08_N&Kb.HE
G(I2b5AbYJX+G<47_g\>K<(eA8MRQ+Bg^.+0PgGW1B#?<OK<b]AHL&9a&3Jcf4##
aR4-AbHP2T58OO&9:R]\CRC@:C26LfK1@T-_bT1O^3fRUHJ1/#_ZP/EP]=V\G#>]
)H4^N#fVRa07>V4DXPgd=(,<8CU\-X3&B/TGAJ^LF]a1C/LKXILRNGc=I-V\X=,-
cTaAPJ=f=\;8W]?5^]+(/@HD&@]3[cS3^;Z,Qb[11>(F\e\bZNg+RH7b]Q)Ja)@+
5Va(>R7F2&&K5&\4P(T^a38e>U^K6=TZ_,./Q654UNcgdT?5(\_CIFY9ZE9.,=LC
#B5[e,JPE.]2V@JFTf4^H\]I[,Q=YOUA7a92I(0,)Ya?7ggGN)?d>/)1=6V?#&.0
Q0TaR>1VB8R8JR[Z&B-PbT-e/RGc/G1N=b#M4&63VLPeOC;dV&IFR.(L_]9Zd6Q=
fdcSdAC&,Z0dg1cT>56Y@J1O0]_BZ((@EN(][>CeY7</1L2RJEe=@]4L)Q,R@#?S
)c95N](?fYHEFW?7/C@+A[E6Vc2Y0dNaGY:_Ae(LS1]dA1+0Ra?:FV]&DRg81VS9
(O)\(9AKN#0J4?&bJ;->^,R\F9&YKH0R/3T,M)BB295E]@8eBY>C&a(eg^3QI.[L
)bF.^0Sa874)99H90K+^e(LQ8]GCH=8?^E3=,8g^77OeK;Ea=,\KcBOXWRA&28^@
1Of5+^59Hf-E^L(HaB2[9JUE3</;bLL8\AabSZKY+,O:<]<&;YZUYUd6;\[5QE##
<_].)e)Jf]K;f:R9.ReK,,O:6Z/F0dTO-Hga\ZP+[_8MW/0JK\7g.gW9STFMEa4a
4+T>7EK<+CYOBNU4-_;FN_N:cNQ,RV(U6&74I12\U8gNJ+@EfG;^YF33&_dE.LdW
44Y9EW;0H9D_KO0H;e=Ve&?+]F+Ae58KT+BfGJV),&SQ,U::(;C&M5]_F@\F>:Y@
+Gd)IQ?DU=c^/O:&W)TSWeME9.>bN?4a=SaWP>(>)/BM\_NV36^D>B[^]KXbX>?S
>6g>&U5W>E+LO,9[^]Q96;[9Z)LEJ:\U9R@MY6A(,(7EX07<_(:^;cG1^-0YI/+P
01LAfYBcERN)@c44:aA#b,ZA[ADG5N&\Y6X)5[,/P#&U^c;fA:G2TJ58:1g.9WVS
?&&X/I6)ME/T3VJ;R(gYJP3=3).69I-\<K1JBINgg/]TR;A39fY>]L;@#&JcA./G
7E8BEURSYHUdZM\4^0Q@0f\M+KA4&9^)-7+Bd1SeVF.7:Ga:a4QgFR?#:O0P/Y#A
RG\0@4UG]V;-D1K1JF]FgO1,SWE;ZESe<=@)aRVO14D16PYeEH#N?(-:S4R9\/e#
&_T5=N0fE<BVLUAQ?DWIMU]1Ae<ESQKKeb,dM3c]6Xf[RP8/&=ebDe]cf_,3ZXf4
#:c1)gVRAgIV9Y[GS0#98K\M2BHWF<Q^\.UMAGgGUUTBW0e+C:R1T#a)SOIGWUSQ
33>MWZXe)(.TJT5C42OKWT#UD^Y3eX:G?&1e&LC):X286MD[5&/VV1/gJ3PU+SY>
=H36ggA>1Bf)D1-STHg+Y\O)\Hc?8=KEAc[B1e-3Dd(WXP:-M;_6)>MXJ1.B#-H3
FWZ/(MMcfYeO.#Mc4H?0&9A_=,/]B+A&(ZB);Gc=))2SIeR(]#?V=YQZ&TZAY_L&
A3]4XNb3)?,JKRG/,8F=C/@<Q&;Mg[4KC?a-f&ZLOKA2@2Sd]0[f+L[g/JR/C,bY
[PG5=,J&6_d?@6)Nb<078O]0=/0YD+QAb.b4:G+F^)(_c4\6L8UcMLbH&^MYUMce
;>E(H0NY:4BIeH@aJ&V_SbBIW[S9IWPfETM_bQ)_gL5(4:95?:<0cTJ/geRU]Cd-
^\If-_+fNL2f3TgV>6F_fEVEB1A]:<cMZ)@#?8fQ64C;Q2X<AX9@c@P92\M+B3_=
D\6Y]UZ\+TaD.bKgGAAeATLQZb._agMf]_21/NYf0,HLfVLGca#YbQHEM.H11.,.
/Q\<XB6Iab,-&+,:S@-acU,1-S]3/cDT@ECfLHHS7M&&)G4(6;ZfVNYQT-P#a5Q=
#RAX_QG2\;O>+>YDf0:NGHRW]c7>V)1-C=HOTNdXGFZ>[d1Xf(PB3CcIU_J54+BQ
CGIc.:5B/>+e)IE,0Z77D?(cT)DZef8[4S?K?9_6-HMK\56KX/N,<c=-=,Q8O_GF
HgC^7(CF+#KK.Ub7;_R:PV>P8;&8=:MV4;:XQ0g_;4Ec=,5YUZAHC88I@(SHBH4a
+V#.X1;?U1K)\bHFaT^U]bW_.GL6SY87R6[K]:[>/YdRc+PcI7[_<_H4EdM>_FVg
<I1T1F&@D,JF=6VP@[&D-+_G[LM6U=98<X)X(gQ+d4KT/aZ8+X;b]A9]BS]0A+HG
]^]TR=FTYT^#IW?W+4[+(/V\BB=ef.)767.P0+/eICND1JKVFNCAZC:Tf9gbM1@W
1?SQZ1d@[[b_V]f+F08VOf=S-VM+U?:NMYH]73_K.@)R#\I0+77RN5J=W(\S8ZC^
K4C&JOVQLKVZGZg1Yg\5?CKTJ:^=e&FZZ;#O>+bdfAK.JEC[0<[K7[-=VUK:Hf>X
(ZPfXeD6GYaM:<ZB:3WI7+C]B_A]We43dBdgN9W9F=&EJ&L-R_Q^&)3I.LTP=YeR
eYGPYT[;.7,fU3U11RT^21LZ5d<9\Ba<>dH_(K#cTE\cLGc9@3#T+4[-Rb\N^QYa
KfFf<(?=NKXa:NT&K<&X[R.G(?._W1]#7G6gD@2R22,DG0^Rg?6@T67V2fGCO)@<
^^IV<1>SeWF3;[5GA@IbTT5-A2,6,83;e;SdMf5;Z&/8@[,[YBgO(05N2O-=dT#Q
G/_U1<;CUY=B_Df#?^4FB5ACd3d+X;<M/>-7)AJA(RfM3L8M1ZC\,&3[6(EHD)^U
>DZR(65M<96YPVL>2C,bB=5:J6)8U&9-5e4E55_HJ\40P?fQ2\(:Q:[&\EGR:M_O
[4@&P98U682+]+,>5/cE4/=&Ef=/W8^BV\]MWJc06110f<BQ5^C&]f[OA@@L6Y.Y
d6,J#B#:@.Z^8>)[^A\(GC3A,#2B]U@c#5IY^1Ea6b)QVRSdageHa>)N3G8<2)?;
YC[5:M.G-LCE[C6^CKV3d1aTFf.;>2>C#0+d-G&EE&O@?6?K^?S_afF1]\C?B_C_
Q1,Md5@-1ef&^bVS?e)5+2FgZ/E^C4EN)<>2>OYYg;/1:e;QRPZ1cZ5;F#;YHAM^
Y0RCK5?S)>1,O-)PbXF+,M^QA9872c:a#T>N],Of@g#)]/]>&c#FI+L^XL=/B3K8
g+)WJeJaZ2()8Y)Gbd/TA)XA?6,++;<RY(>N/]BHPW4eSW#9=Y]9\#STUdbO<8+d
2ERd[Y_Ce>S?BAGTLbCQS(=WC,51OKDcY&.Lb6Q.ba\Q+4Kb@S<B\BS2<CJXeAaX
]@aN6+1W/;Ec/=M+[BI9SSF(PKE,Y@1cgV0HI]eTMIF;19a#L;d4NJ0cP=cS1O5=
35KS>4GeTVP@IQ;,LH4QZ&Tb#1g+O,4bXXWU5f(1(7-YI?cMK)TED>?+VIQeU;4?
Y9O)YT1dOQE?FLZg)S[\QN4IY;3=;,aG_A@NP,^/<7#7\>EOC8DfWQHX)@M:N\.Z
=41c&>fBLQbX(O=fcK<8+8152V=&S8G+O?3I4eHH1.=5_P\Oa8M4Q+M+cKB=Nb43
c:W)bX(OXff07AFIT4X2]S]=WR^^W)P8bcS)&>QAe+-Z&<:WCM@CP[ID8.CNHZ/G
/d\]-YP_^a-Q+QSYbXZI-WaR=D60f1-A<VMf<R;U=9SY/;CRHB7P.O\5g.UZL_DJ
S,V)6M@F)55g=#W8/;1GaK(:E(LS1Qg3P/#PNfgN-gA,Y0=6.Qd-c)1e@dU;a--9
G@S:YF);(GL21S&DE@M3gWS].7G<(CCG-5/7UaAJ6K&6g??W<#^@)?e_@&[-.aB]
E)6OH@MXfeMH,=WHRgR^>T\@A\Sg/21&VMY+ELGV[eMgSS+@/adc]Zf6]NH@WU4B
NTH:U(6f8QdgK).7?gF6_?UC]adc8E/RULYFJ@gY;VXX?KEO]KYZZbDT\AW-R:<H
S<6,f58#S.c^dXBD6GQA_+L=#4PMFLFB[(C@)f;/KNf^]:,HNP&b=g32H8I-_8=4
]]N<_(V[_MN<GIH>Yd7;IS>[Sc]N5a?38,368SGcP]e0CR/W+U-:G]H;1>(LKe(_
))[T;F+g)-eK(Rg&cZ&f)TaA@KZY18&[9)6)daTcIM.M>BMS1FbBb4L:WTPKZ?9C
=7.<cQ39P0-I9X11\U?F:SL8LNQ7U&/43,f>cIY#Pd2-^(Tg<eTMD<6\>aeg-\)/
Ea6GW@a0eUbZR306&1#Ag5bd+=XD&Z_OdK@\,Ee8L^LVKXG?^:FfFegNZ,-(=]H9
7#[?V&5[aI00+b5:A(5X(Q9R@Q[#4&CE(ZIf7dK1&KIY\N=aFJ0HBD?\VPM]TgOW
a+.F6A5]BN84cV8PS(B:cDL+d&L(UQHH\MbZD8J(C#f=fV+]=,g;NR5?G/;DJ?b;
(/:M]L>]&,F&Y03K42;f@Ye/?^;X@<6Q/<W0^6.(&88R6e+eFCRI^b9/N5gAWRU7
(N0M(cg^5+L&gXJ4KD-6ED35YA4.QbeMA9,)RPKFK,a>\XC/dP-JUVKT[.M\0C4&
KRX<0-3]2aH,SA/C,gZH+B5L\6O;TN8,N(fc(BATGb:dGdCT2-bWGAJQ5P0ZN77>
C2U<S#d6dEWE_DL]C//AVbL8/X<9PEX<#WH5]Ag@Xd?db7?4b,\>GId+d4YbGW16
90K95VfK63?f@1L93;Dda]#246TFM+PSF9)F&If\@gEd)C37\5G>3c.IAc2[_,5g
JN]V3:NJ/Hf^_09HZ9>e:.<?MG8G7Y#0B&d\6_+]:MT6;W7WWMQ7E62+.B,c2L](
cLT;g>1O+a\ZONR-U<SVb9?13O+N<aXO]gLQSS3F&U98B76JP7>1;PL&a@K:492D
Bf/@dEZ.TU<dJMa@P^PbTZ>G]X3UK,GIL5RTR#YM@R?=f;3=]49RI]P@>9Q-I&SQ
4]X9^P0VO05((S0)<#B\_SPP7PG\8;Q=[c/MFWI,a2^Q;74,P4&RN:@OWOb?5\2C
50Rb]c=+c3PRWK.)Hg=ZRdW__S[.25c1:ZR)&,\?J(4g+AVfLf]@BP<64-W.BJML
N@-K7Rc]Ic[6f9gdMVQbE^4,VF1@CMR=_(@EIRB]SU(HL@M/Z>]e,BN2B?AO6B.I
a85dZHH?JT1Lab8C1DW<PE>R1(M5N0B^B^,c?_g9bXM/0)>I(c;&PT+R_bFJ]VbF
BDQQ][)5UJU;3fW][-=:06@KQ:G&HVc&-29RGUQ@_OJ@U:(4#2d5VL;1>XA&J).Y
.XMUDO9]=)5:eD;BRa6X.3CN\XCP\-)WbZ&f[_99S.>=1@e#BOceKL-\=&B0W#A-
RNV.)bK,AdGT6MYSg+L^4>0D@RgOQ[eQ,BWPCE@48VET@>K:@\2_(NYS7X_B;+:d
_R)47EYKF3^&2\)Z<Y#@<S:BIHZ>;#IOE)K<]f2\JWN=+W5+DbU1.Qa.WG[FdSK]
FN5:+=4\2ZD2gJX3@?Ff025,f8T&3&1W.[Q,M#MR\\cAcI<EKTG/N]c1(,>)Td[E
d4-:cODZVV<MO-,2HJSK27:(=5X&930TXR=/:,#T))9^=2.A]JRIe95&MGUXL=<8
#(cA&]M7GcDK&^=ZH1C>[fQ/LG-J(8ege<KcY_>WK^379_ZSF-<3Q@e4YA]=LcI&
[)@O-SXd.J7@SAOM4,c#+2=Y(DQTSP<H.NP#C6eVZS;7Rc,.):.8cWKQeY-@JW:.
7V=Ug;-3V&4,a8A9a=e3gZg9c0&P1K+J6VeR5.VU2Jc#.[c0c&f<MO#3WQcXP:M-
78OTVPT?LbP32>MB96S8Y,TcZVgfO,,;IT.T7fEN4^L>b58M2;Cg(Y=KB7:H-G=H
0:\]0ZZ6?:XJ_X?Q+),TW#_5f76R9)BFC3_Xf;T:L7TG+C4e0Qd+U9/=&@&UBMV1
NEYQd#YD)2OTX#UC.U:ZCd8eI)(ZM,2/A93YM.f(-UNR_D,)dRPbe8SJZKPM^YG-
BQ,f4W4(b]D#Pf8LeVQDV;V68T;&CIU<He#@QEY)^01T)A]NSPK\TZTf,JZLdd#:
_=a.^_^7b3?V_L3J4J\I7c)9STd5[X#V_,UM3,I>F9^Vb]::9FT^J1d+_<Mg-J,K
#PE5DJ;eg<KEU,EO&]#DT]]?9f&6f^^+/e/\Q?3#Y>fe+_4\].B>6UF?&3gVaG.C
O?S3/^Ha<Z(3>VH+\JaB\\ge?]//c7RR9e_+:>K3@L^C+XND[/gLbSE7?a,ULY@d
B>U/BF9EO4QFUX1;BHK7R(S[9\84Kefg9^L[3);U>R(A8=9://3Q.5V[W:P3Zf@O
0VI-.FQ2)3d/DDAFR&<KO0?1Gf(.,XeRH=B+(f#G9X[^_[6]bK\)5-,==_^^W2/B
c25)ZK&K@XF.106I:WE?bR,I:2F9837(GJ:cO[\bd#)Q^W+15I8N@;/Q-4U@&P;J
+c9:[KcU34CMWJIc>EeP^\HJ?SCQQ<QH&-B.f94A5gES_AW4:XE?]S;:Qe8G[:b.
1QK>=0I1WL4IR9N<A&0B-10E99d/R);5?V5=FNCV4(^8W&,7@2:^FC99QPe@24c:
_WEDRN3f9b?D8SX>JT5999a&T]86;cE06\[<&8[e>4H79N;?f-35LI[ZW5PH\4BE
8_F)caAINY90R2ICg.(V@-)9K+AE^^57RYR8?EX)FX2VJQc6QD]A@=<0B@GMBe\<
,37LWO?Rb(ZD:6#M;&8_H5.FIY[CK<00aT]?<X?Z.TL9+R&NNY=;3L?(d?ACC598
OK8V)P0..91F+MH-\JBB<6>]T1-Qc5S;1IQd1&X\/PLdYUV2d]GM)b]6ZGfNJ:C2
_77#dT:::R_[7-[Z+-D:cOOUgV<cU:94.[?,X<JV054cg&0.YUYg^8FO[5dG&G5C
^,/NYQf_=L5NE&ML-<@NgaM[gO5<PYbb(T>-Y1D/5,eP-/(09-#O/M&9R6]8cB8@
^/^\V]>+A;#,AY\cHH(AaY\Kde^<.QK4HVM058C8Q=GM0DWgX0Q1RA>2AK/DSUZ5
7P2]?--1Vf7[=&W\L1)XJEC&+=S]3(FEf,5_#fc^aKU76CB]cO&Q4_W/53;Ha<,M
Lfg37NcO1PLUf/)M[eSF._V6C/LQFUW)/G[-0HA^ZF:)U9\U<\W)9#ZIdV;0>)BG
VGL+^\K7+<NMA&H+O^\g@a<5=8C:bQN.=CJEVQ).BA_?E7HLGg0#VXN5b3]RU1_@
D15O7gU4O^d]5VTLSZ&_17V8J9+3OWa\8EA1&FXKafMTA,;W<cTLQ^Ig_G9egM)R
a4UaNNgIQ>8SC+HNES+P3b:0-I@,^f>^]WU>MQSQ7JSM>dTO8Q@fW/b00,IVAH,A
NSXY-352ZfH7:8V<@1,fCDX8WU:ARA4beE<-Xg(R62T?CESf[-RC&dQW^;--2[\6
=SEO\;Jd+0Tdf+QLa\GGaXIbY<B;OfRR1)gcB5M7UfGKW&c4b3.aW#(F2)]^VS)^
J.03XVb7OQEI(e)[bcR7K],0D@NX;[7QS[U.3RO6gO68FVbS@3-VbNTKO[H<>Q+R
S.ELD6JEcaY+D7EQGBC=bJUAb(Pg;/=UKf>_19+CE+]XM/(9+Z;.;S@<B:5.8()#
GI/gd2C3;f-FZc158.15(eME5Lg5SI#K0G=;R/f\S4KU)eAE1S:Xc[KHa20G]Q]8
5WH-T4=4V8GQN1DI[6>:8&QZP-4Y)=49K9:\+13C\(MUdK2Q21a=60C;F+89(;0^
?6@cTJ4];QWO?7g_@d;W/ZG.7:13e\>(R\b/5VL:O=S><9[6C392+OE4V:7dQB1U
;GQKRS5Lc(2#07NC0F.&@;A^d>IS8(/+76@R8UL+g_APfFcRKa2#+cgJbT@S+S-Q
J_B-I49_SY-P++>/eRf]9B2A1g&bEWBPf-?97G(VRUH9g(RW?QEULL>]gT_c:/KY
YGS^_G2/I>/#@A0+<RD9;8ZM5_eEL6a-K04P;VGJLJQ7188f)F72090DaB?ZS>44
YSKcG439LZ\1_TN8<+\PJLWD/=_41)39,M947\+g_GNR:[\.J5@-&B\ZV@-9@eSC
7a6c6^/>WR3]VDJZg#E)TgMM:8:E/g=aMPAWUW-GIOFMb@Ad5\RR(Y68-4@CZLec
)E?eC??LW#LOV)a7Q<S+Ta&N^B>)67W@(Ib&930&8)0MDM47&P)U6FVaOKE^=SeM
P1#)BLTZ_J4Qa8PFEW,5-:d9V0EeEPO;/[N+I5;6Z7&E2^I5H/c7BBC77+M(9N<P
<YBed_^0Q@;@\V-&g4.G;SRDdF/U<_9W3?D4MV9P@ab;-4^R=X+egN:\)QS^5f4/
CZc5Z:\dW;\T?;2dY?aC+6,#>NOOS-cZG83dQMON\f>8U+Z7b2,ce^(MND:9?I0V
R0E#g<V)6aAaaRfg[A,+\D\MZLT#;;C)@?[aPHbaCU;XEE8fYNIQb3O[C7XKGee8
TIU?06ZSbbKg<_4OMF[4Dd0QLe),PK\eL2H)6gfB,Y+Q507eI[caQS8C[P\<JUQL
_7\Zc<0(VBIAE_[9<05ANg1d/3g;61KO[bd)OELKXLR;IGAIVZ<\+EA_#O6f=M-c
25)68LEJ2@FfgY1RM)9XMJe8fK/RZ?WIZ^0;V=R(93b>_2Zg-dSMf#\ENSA_][^(
J>7OSA\A^]WQ)[bH)#SVa#V[(.1+D-G/,WAd_\^a.KU<QOf2T/AL7.6bSfY\\PWJ
e@EQUg/G2X[)F(<g+K8Sg&VRF6427W0/(72Fe@ATO9b#UE,<YK=fc2bV>B7D//4H
.-\EH[1c\_?(1P]:Mb+X^#QU)A5^]\IE_Eg9g08P:F@7ca6K(dd=?>G;+Z]BX+.O
H[(D4Ya2&>:O[0dBH-@KV>K&ZZ=WMD2S06X[EPI,HO1E_:3U3Y+MBML\LGK@5GN2
>E)/2R6:Z)\M_KIOA,Ye:D5]CEE]/6+6()-aT-\LcL6WC1UAZFJ;c@CCOO\U>P3(
1[NQgY#6EEd9(:;O<_-G#bHM_ZF[H-;B^.VO/>Z^<0NVg9(6=J)P]HV-P,BSIPX7
M-7FT4b@aS/V3KPHQ/U-F-91F:C:bTR]X,E62IUSF.Aa=^9;S\aF3]7ccXJeZ7NP
XXM_OB#_._)Y(@Ca:gH=fF9O53VR:e[8/>2=UCQ_QF&0#:N6GaYI;QDUeMIgVQF7
>B&=ROT1LD2FJcU7LRePGaG]OONV05fC:\KAHGc>#_D43ZIbX>,TR;=3C5UF_)aG
e/S[CI(O/GQAQK)6X+H-/9EV:feBf/7ECR#7_:PS?EMGN8]UVf8dH;GRH[-;8](]
89-8QKBTC&)9bKZb-MN>XJ(=_QO>M)^6bDX\&HEZU/]G>?bZ6cf?4:FX6#NGPd=:
;.#OMXRURN)==EV+]-IU6=T5E6]bW:P,b^7S:@_G>)gKbV;VFM,ZCTC)Q@(].^D?
Y[O^307)a&D\>gGHfH-<PUaH/P#D(?S;/Eb7#&-;K/(U7aH_D+OG6SW06U+YSYUF
a;e_0^9Q,5AR)&[&I;^R+6.K(+HN[7f&60-cZI+:J<f,60)aS:=S-3Fg.Mg_<MGg
@;#FYLfU14^V4VWNB&S@(XE3Q//@c/@F-H9O@B<+KOYCSI]FGD]V(<]1aKZQ&ERV
K5\\\+K3Nd-WTGK9Egbd2#L:OYELI9ZbT2O/9:dM7VeANRePeR-PRH2dB[5,^Y)J
W<Qa8QZ+GNNEBg;MN,;ORa@#?F#Zd5]::-[B5<AKRCD5N(<EENA-5@Z(YHc:_KU[
5U:NJ3\7\QX75]KE3RaK#A3b/+E57QA4+&Q7fFff6IB/[F9(>8/.<O4OL.Q7e2Y&
#dW3b3e9RT?6dNT(;dfWegQ(YJHDdf?DW&_g0C^g1H[?P(2=UgJF7EdQW_K-VMag
OG1E+B/+F6?^)Z6-Q?OI]Z\#4SZRd:>9W&cK=;5(]Y_T>\fgJ;U9S=gPI-90X9G7
:FOgD1E]:^&(a9T1QD&IOfU^LUG2a;SXB>9gJ2)QX.(3adf:a_4\_UR-NE00e7W;
XCS.d#^E)g^S>VP.&7JN\]D561+?gGT\MK>^BB1=@^ME<MW_=1K-X^b^^f.M7LFV
#DGY?TX8PH.U-=(Q=O(D,>J13d?TgC/WCfYOa>P7c20d@S]+Q/,/fIP(R(&0+GBX
SZ5K&eYJM3>4A-;YdCa4LI5A\53+V3HT1Q6R,G,gY5M]\ff[A=f?99S.>M(3A2VP
YDFf7-MKM10aBOV-,EA<WQcZ.\]VHL3M[[Y?O]-a#+=BJeE<c]-J-/+GeC2E\cB+
5E]@3H_XcX6T@?:8&bPO>2Aa^c&D-)0c0_=gF.UAf<=]3_8)a;5CW,0/#G^fc17<
W4He,_AUNT&>1JNJ73/aYFO?[/c&FTRg<0JOa)^A.3eIb-,<I7X.QG6S=KO2Ma^S
b:b<0]FAHeZGg@T-C]H@-H0c>N.:RdQ9F]I9Q(]S+I__2f)a9_3ZW:O5-]\1PQ;J
9S-,R4F-(7E__,X9(e/aD.6&00FcK/YZIX6f7OIX<_2<UGA;OUXcZc\RM1d)WWB\
e2f+Y[_:6JcUJ642;[K3GT_S<Y_/J=DPbd&0TF#ed^0Y=65N&3ZRK[_[G]5FGF#I
1:B-XDM<T/0Uf??>Y4ddfOI\d/.TbcB:4C-74(HL6UZ&:YZ84T?Cf8^Zd9_:E.BI
\IXH27)MC<V0]//#3_5We2?X3f7JG-YIe;NDgAFbM#+gG44\P&#]3=-O.E+D)HfH
=PVZYSKcM2O;89]BWaU[AZ590R)\5=1.?^9UTa/Y_MEM><-Na3.42ES2/S)I;Wc@
+@XG7NcPU2S3aD)@SXZ8DYKGEGK._ZY28(^JTGR9Sg<^^;RdFS,(LGKFOefe@9E[
J3Ja]H=A]/Sb/L+QZ&K16FZ.KaTI7.)&1C&US9b#>B9(STTc[@RQN8/ITe:Jc.Gb
E9Q0fGRBXO#Fd-W?[]T]2T&e.aB<J107]#Rf=4g:f7^gOfcV<MFJQ(A^D[HMCE,F
#EZYe.\8Gd,R[:PA[KBE3ENL^8&4.2HNLQ_&=Z=@A@3&3E6P)GB52I65gXRbb.G@
N1DRL^.25+PDWZ[JC_-S9M_/_FCNYL8f9L/Y<a44;=XV+ZLLA=-OBb?_JUA&e4FO
_+CZ;G?MQ(LYF,4CR^@;F?T^+]A]4&eKbEKe/Jg4;HP-&D7E.g#H6W\P5/7[2_@E
KQa055)C-#JE87G8[gBc-egGO).#@>IDgSPbWXISdZ,X]OWb.]_?&aUOY?2PKVTB
a)LX@2E_P5.?8P@LA,\X?ZK^5e+[8H5M4RA[PKF]@]a=(0A;,7D2Jd4=48d[H10g
&e.RAB57;<bBWJ):JgQ(/W&H1OQ\0g(Y9\O#U-Y+EgWc6Zca2K9_L.P=Y]abCV7L
dWV.V/@&9::X9=(6[8U&&1A9cBF71]9e]gJfAVAI;PQFXT&(c@-,eGS#I[/7WI_+
POg,dA9]eC][W=/BRYS]a-K96;\P.1KPfA;)B^QbHTEfPHR8I<46Wa[eOa0V>@?e
C>]R++7,)B<@B-aV844e#-IS-2e-:KOY5QGg35.YXf[7CU;<S(9^D+S)cA#N#UG.
L8M\5G--+E)g4OZ=S>L?2EDS\9g-,IZg[F#/BWB/K8dT=g_,;<gSQD]7EK&fUT^V
T53?UQ3RPdQ/3=/8D+V7X2NP8BN].A[6Z/IW[<8GMD1V0A8.,G0\LEI@AM4P>NJK
d]OWJ16B^;=/FR^/&dDY@KO9RC,85BMEaN,X-c>])F_Fe(.IVF(=6c].G@B0YEV5
:8EH6;R?R4&@ebURV2>fMT-1^I6BNIMT2b4R9TSf>6^PFM[RNa2<S#D0^@0F3PP6
bU.D<X1/^?+PF&=K@cKUZG]DA:M4M4g--,COB^,57.FG40N1]NgO.71@H.8A&b0S
9LE\4[CC]1a^aKQ.L?]LcRWOF99ge<RbA(CIOLJea4M1SED.,K6E1F;6aFZP8TMJ
U/9<LR.^D2D_1TX3J-bH&a,1)G-_RZa;f\R?2cFSOX,bH+[fU/KEKMQ^^QN3gT25
#FLeW4U=I0QeSPBKVP96+3W-#I>6.EH;e<4(LL#&CC[S]V[[/Z^2g;6XV&MSU<gf
T83.L(ZA@9+]c/C&KLdHe,G8.GOTa+D5(5_B+M_(T]Y>+YS=8E^NKYQQ=L5de:(>
3JI8#ScEWI_g\+63+)90@9:a2H724F)7>c;W)WPM^.W>HNXf_Q;BCKFHU#>CG9E1
155Y:VXg)(B9XF-P<,A_e,gae2Y6.C:,<ONGa3?DT=Sfb4A<(+DddL]a>G]<I)b[
8G25>UDdbVG5I?SX/Sd[UE9QaEZ?eS:PGR.G(?/^/J3^.(_81/<gOPHP?7:_9EZ[
[8\H4)5Z(AEM=KCE>F[<&Jc4WJXfMJ3:e3,A:H/#?YR4\-EBK7BOK)Q=D,[NT=:N
O/d/eS-O,.T\/)1f;:5&7WL&bUPVZ0)2#K1.6.UDeddEZ0XZX3((B#cILeA>3C1+
D+D23XT)D+MF-?BeFM?=1SQ\TPFAD-]b17RaU:K=P>.6#-N2cHM7[db.@Zc[UYOX
_(-O/R/d\AI0]cYNB&Ea+)6/^WBB4QEe7Rd:(XM5_[OUQ=PHfA4421KYP(7O0Q(,
4II2B<#)L6+Y9EYLbV58_/=+?F<<I/U];R:G0bU(H;E_\TWZH2W[dV<D7cBF/7;?
X8@Y=LW>G69U1c.b_7Hf)GNC^YONZ3VTHU>9_^g\_[P:Ma,D/M_.BQEdV^@:gD=B
.A0_SI]dE;/N_\3F;>/I^D4)5@Z)UA5UaEH:L-H<)T>d3BXC6-)TKIOCa7,b0c6M
1Wg.#Dd#e3M&8cQJO;K4SB-aOffIO^_LF,d:1+CW:BISd:dWK#E5)]<EEXD;B&E9
>JL,e9[RT,N&VSE^fPf3/BV@M>[(OBU.V+SZ0:QW-A/bJ_g.Qb#GZbAV11YSOJQI
3MH)F]C:)P\VGRR-UC&=5SR\W81T;Fd>HUE[:d,YTd>,_)KVWfY4fT;Qd3<]bIF+
gN]d,O\0-D]NJ#\9L&^R/0FR^c&d:F]NK_f[UW;)MU/6C-,1C]4/dZ@gDK?#/-)[
84]60Z/Md/>C0/F[6<>:VJAe^-H.WI[N_^3#==;10^aBSA6[3eJQQa;IeIG6Gg.)
6;6gPP9c>=/aAX\KD#([?<-fY+XPWXQBe:YFIAI-R_I/HdYg(g+@]AFN@(2;1_EB
#5g<c_C-CPFIA.1-CN2dHZ,-O-:fMF<.HbMXAHJb@aJObL>MMYH;D#Z77#DfGXPZ
(Q:;,JF;@bNDHWIFBWd<OaZK#4gXB-Ed86>[6eP;;_1=A8/,:[ZMX@E#VdCT2WW7
f?3[NI#RW>2SNMJf-+2HeR6,+HQS)12EPAM>4B[aK]T>g@>=/0C?4IMRMF@27/2g
JNKS&AVYcf=&^@f25a;g4@=2S4C.VZ5&,+7ORIT^M6(AI,A1d[ZW-d?]?]+Y9@MI
^UQZB&OO@d)d?=?XB2VI8=&&)J;.9^IK;C&bR^<VMZUPf-FYRd\a1c<T@NF59JX[
@CT=L2M3f</LKZ-FY_OW][a/W\S\->G)()AT?ABGe(E>eHfUSeXd2@f<FSUD0N+W
0ecJfL0&4GY+X]dR.-A6OPU9Ue(7-IKY/2c7&caX_=PM0#Wc[2]LHaHJ^7(P;0=I
[cO>U#&XM?777]g6#?DdY\8@JgZVDQQP-=a,3M?85@/LYIcaLK^Je]dT/DE(bdR/
,>WKNQXD0gIJ:B5eSPF;cfWNA-/UbT8H3^1R>Pg0E4=QBGR\??:ge(,07G(E[U>-
e32^?/EKS[U-30^&+[)XZ8H]0?IU.X+D7fb:d1)1>_P,f,>cU0BL\T,3^M-S4A>b
f]Q\6=?OM8K?Eb\>5W;TGHSF4X25T3#5/2GBc-@NgO</([B?[CLZM@9S6VK@gX.D
]abS1G+B71deNXF&?M0.HVeG-0[b;60IO+0=)Z^P,,eHO7NO.1OQBOB3:;ITJR(:
I7.4gKcAf7F,#cbddIcK\Og(:VFBEc0f=:,E5L>()&Mf&;Ra<>fM=SIaU?;O\J=f
/_4]Mg9fMe,#fABXd2C\,F4e<SGU54L&-,.9[C?BY(DA:@C&YCXbXLbaYBDX_-JM
4c5b9_f/PK?eP=YNTEXc]MWV-b,1bE1&T-\ZDB>WW9(eOC0g0^[D#,JT,;V=)/[N
F>b6(cS0BKcWU;SGF=<7C_dgU4Tdc34b<D0]S2VdEVa]c2gF2a#G6B>E/]8]#O_T
0,/cgS1,;Pe<CY9.GcLM=0?^Q9BKe]]WDadZLA8cMZ;K+=MI0C14?5#=&@Ce&=>F
fV2-Y<KO\ag4\J2aC^QcA<Lbe)M<]c;7,/NGg/MQB7e+]:-]a6g3;(3-OGdag3c8
3TT<U_L-G@LeY:Q9b+@@FHQfPDR2@/I8L.5M9N2.\IMR2O\1:/-.5OSfMRA)eM-R
0eQa]M;=^RZ&HWcJU#5E>V6V=+1ZZT+a_76R#J758[>P;8a8Ffa,\@B5e##E.EMI
-XeUG:OY^aP:-[EO&[,0=d=08CF4OeA9aRKR#T](C@ML9?S6^5-8:WOGX?\=YY(U
IUa/G;e\e(NQVe5+G_Cf&E5A9A:4E(L6\Yg.9^/NYg,gLJ1c.d.X-#e^:^\_7S1Q
+/PS<JNPWB3;\HVb^UgPT<C]O+Y>GeNZc]]TL&]#d69AQ^=B33^1F4Y0&&QgI#8C
a(07\bQX(I5YS]DGaE;ISS;3#346)&gH&_@PC@UEGWAVac\f,OAea]Ue>Y.B0GDU
#HeU>B<)fbge9J<WS^>fDB<Ud^O6G[K#b4:4T6Rb+>(WK1QHMM6WTLLf-M)#==F@
5;HfG=?&:9,KN>c=fM)F45CIVHW1AU,VS,aebA(^O_?-/)D2Ee<?H,>L)1MX3\dA
(eCAaK>L<WEW)9G&MfP5>;8OcLM336NIWeP+d8_M)b(E#CaW+IF?T<:#)AMXQ55T
dG@+QH\?)MXN,a.02/<TNPI_1?X@B5(bLN7a7CX:^<S8aQd92)3/@Y]E?TN1,9g)
D\>L_Ba--,N^\-bLQ>fR[?JK&0g/P;c2;=+C]A8Nd&=HRIU=/Sa&>TU@Y,A/7dLS
B9,Y[5TRXHVV7LWbO4[VVQ-<4,,DT?Jc(4RecRBaJ8.cXN)YG+KeeeZDD&:,@=Ga
=JQ/0Vg+CKbY<N9F[>C,S#;#Z5A0e;@M)AXb0_KQ_6FGdPe(L<RN3WQDe=:A,_VK
Pf.B=(4ST2#H&2J;^O>ZICIB.U+@Cag)#]6.?b,PRL1&@GcdEM#POJ=HeL;&O&E<
EP2D9Rc0YVa#dC(bSDWGS\522V>a[E0VJAM?CH?B)2Z#a=_W][8A;XZ.A<8R\8C2
[B:_I#d3VCFb+G.[3+L20;;Y_67GdRd_2R5O8ZO6QUZ[(K<R-aH\9NY?ZZS]J/4V
ZCSSO@<&#HOd^>Z/6V@CI-Hc28^#P8HM\g=QM@Fa:9:B9[f_:G]K/:++OKE7fTg6
#6LePS>+H1<Tf(f1_60Ff+(_c78JgGG?2(_.#HQL\&aYWa.X?IZ-b?I3S:@C<M^7
g1.^d8)K?&_@,V,OJ4J:+eEg9&7A_9Wc./[9g&3Y;M/30gOFBM:a_MCLe:baVMaI
&=[9\4D?[F5:PgdF;5#[^UBdP7#4[gJGB>XcY5FVY+BHDf)6G\8O,/4-MGRJ6>57
e4?7XAXB@GC/.f5K-CIeV5E9b.\+5,Ge\)g,Ld,<::f.9UI_GQgS,#eC(CcZ^UN^
Jf?)BZ,V.YQIL2]O6EVg@W6a_TcWL11+g(PVE]Fc5ZVTQ,/&0RITC.Eg)Z\>.C42
-FN<fEDf;?(JU1J=&4K?ALBN+<G(-1/G^]MO#GNY/NCC&3gGSa^#SVC\SMfca/I2
d#[_D[O<?S+9VTE6USgKO1<\g0I+2=I,fAB]ADa2CO5;VM;B=ESbZaRBR86=ZRNS
C+I?XHL2A&Ad:U/QUN]/^+F>bIV5[TJQ>UZ+BWAIJ;Q84FIAZF5]C(PfcU1VdS2=
Y5:^AC7:U:AcLW_C5S19fBRU6Xd-A^MFB&1+[a<_+72<[;5(Z88LBMHTR+aF4f#4
>2cc[8R4DP,J;Y^#=1[GP;P^C.9:C@\O/4M82I<8BL.XQN=L(IT[agg,dM_XAG6^
F+aAd=,^FfKHb_HL4SJ@W]3J9/Ra>/.5&WUBSELM.a#<Y_R9-DPV(-]>67Y/5UI5
W?fcW&XcgA7)=I1\/6SL91eO#;?>9&]55-aOgHfM?FeR;RG\UKWTV2(=bYI)F5XQ
_5V-/23dTGGYK0Z58fSXNAB[KBI#[.c6:]/bT&4aC_d0d_HI)-IYB,2]2)b0b=)L
#Yg;R#<)+K5d/RfbgCHe4&c=aJOPTfdEb:>1SJV4]0\Z2ff-)C.Y2[F<,\YeDMZ4
(0b#+6XH1);=MLF[gKe0>PN)(NGJ(-aWLYa29N1TE5ec5A3c\ZQ2#R:(5QDRBS>U
C1\b2;P[J@PVf<be4b,(P);/7SWG,NZ>+S:G;#I>5-9gXL2TeBYLLGHIOW;V?PL9
G.4D:8=>XT678=cQ&O0f];P#CCT19,]:LE,4QMc=[S)cGEc<WV4@d#E\(AL0,2O)
982FGR0gW-)\[W#+);W)9[SaTLcVD-WL@01(HNXU?4QD<U\_gS?L09&<?>]YXNY9
g2OZ2JLfScKGe@3D:2+IeH0_N1B:B2Dd:dQYa9eb=\ZNf>/]<Y>c3bJ6g#@=ga>9
TSB([c<PO11S5ET_Mae;//U+<I8QM\82CTG2RcO,P^.YJ_]Q3NW6+Z=Q53VJUaDQ
_H0I@+-4edPL#+PQ8WfHK>c>T3aNNJX#)]8E&a+11Z3F(/8&#F3.b?>M[9)]H@KI
)RR-)R&INT#g<.Q=0+7dPGB4-EW9,D:1^.47I9Ze?SA;g;DX)5Y#1gG(gf?H)1\O
IR_N2/-9GR=;1KN-M6C06Y_ICU-,N(KL(E;BV^D0=-7)B=8,/d@RJP(YV8W9;-W:
FgW2;aQ42F2,bd?=B\7VY7I7HdHS=34cJ9N-33MD+;E]cMSgHO7,I/((c]QLaS5f
Re56+TC>#SNgZRTOY5M-a1_7Q&TG<HDKF)7ANfg?5gL6(4>HBGK6E>=PLcD,e,@)
B@f#5OX89D-,&QDEC>LE[>Bd-MSZQ<4MI9PB)1F[K7O4.)ZHOY:QRc^F<SAKZM;)
\J1LV;_;55?^XY5@RY4B([J<;R->S5GWX,Yd\RGA^IcY[.XIH,+LV&W1EgZ&,5:\
(^\VE94#cJbEG[L]feP[WVR2H0WJXHaIG\e^\CJ=NIH2+1Da1]IX95KQ1NbNFTf1
_MHGK_5YH2]g\_Ic)5O3((K_AO?56U660,WXKUN8.;GWGPa9[0)aKOSC@X-/_>g\
N>c&eKE7Rd+:]a-C;(TD,Q4B84e9DEKV\=19;/+5XJIN2ZX;)IdD5+7^bZ7FF>8A
<#5.d]NMMUD5,+UO:?4aS+ZONa;b^@F-J?/bU;^ACUOd=5>d5^Sd]4f4BRT2cB1e
8AA5-[F7>XAJgOGcACGCJ/5O]&XD>f(2QL)_E1(C]B0^IM9:CB9?D68Z?(=5L?\3
WfdB:,PNT9XU=X_/=]/.[//O(#@YaPf-^[:;=LP[.LVa1b2@9L\7]M3G8]IKV5M]
).52R&OI+4g:#?Q[b<L1Y&5M<K[R6^XL_A8EVN9A=?[F+dB&eKTb+#Q0N>=PXX=D
GV_H#GB:c,YR1BE2<DO,>/.dMPLN:7PW9Ad\/&+CDCOcO+RUc4f]MXN25WN@?44#
USaA9W@Y5-)VB4M.3N(H(P8NB#Y=/=TP^=J4M[(2&_WUKN\4IJ7=US?gSE/N2;]5
&J)0<,Bff8]OLX=G@<7[TX,J3,K_MQ[44U0<5VK<Jb2MM.B^W\=PJAJ=(4R]2^HQ
B#WcbIC]g&6-+TR..8.gHQY,=IVI5N.RcV;&b/9#):L7@EJR4=T+>dg=/:A:0KX^
C1U8(_e#3@-[-YF86>3S9DAAA:Dg]WLaN9OBTbDV1cT<0WXQ&&GL^2Sg[EZHeJ[.
OCHI:g\IG&UdgDV>?dTf33)]<.-:J_>d,I_gZV[^(>2PdCAb6BTgR\X7]-Zfcc=0
WMR+R?4LC)U<]7)f5/<4;RI23TKJ-?#Y(7K4PSHPLVXI+72H#8,c3]+JSMZGRL65
.Z<XSfPFY2AG]CHLQYJH+7\c@IC_]PSRK?T1,Nbee&b+0WNW6Fe]=LY1Ld?51c1^
+;-:TIQKDZG&8TC(W&0Y7B0T/9Hf#>O=7G#A5ce9B[LOC&Q&Y(L^8B8Ee4QZ\WQa
-cG9A3MfM+8&YHB_L;<_OBdfO/FIZY:P4V_8A#fB&W-KE(8^\EWa_#@OJDR,cRA;
DXLF(:Q9T@(IB7>XS&\a+;FAG#^(+_7)<-/g>AG6g>&AY02HS6J:AB\AL4Od[T^3
=LXI0U<gX0?V>YdC^>BM=cQV+L)-d;^IAD1Pg/@5(&YHIAQPYIUVe50ZM2<:O.g6
1T=3QTV.N]9a<5MO>AC;d-0=8AC(Y2Y\K;HaC+/SMb/D2FX]-TFP/H^.H7[()2=K
[6\f-\;-JE0&ECeRQ\aJ0<V4OXG#H&/d8Y@@ff?;]D01d<#NL&K<G4HL)cU=C8-7
E4SH6>ScQ=^BdTe4#FU1a;ZU/4Je<=O/KDbTZQVbKbVX5R9W<UJPbgAK:d>>MB9f
TYb9&3g.Z8aG0U5HMQ2ME=>1)KC-,b6Ff]728YgZIc]DG&W8I1<>C>N,&W+(/KP&
Ua[RWL<PP6ZE&20a[A##-B<aHG;9eCAKL,UOD3XPAeJYC23e(,CEJ]FaS)]3ZTXQ
1&FIQ^?b<HQN2OB93WP[L_HE1^;@d/+^^TUA2\;-=U<;gM&M?;O0&9+XHV(,WT^>
E[X9g,-dRgX=@T8g8A(6,/_e2@]cE5AJ<=9VN+&a@1PA<M^)Xg,\F_C_MCI)>#P4
NTNKCB;;eUb^M+c87_[g8+[9#?JU0GJ]Vf9NFTZ;-)(IF3<-V.6Q[GC-cbbB.<7P
FK+C0-;XASc+9#G)F3#W#32:(S]6,WB#d?,J#NAJGHRFW:@?IX(._3#Q)U+XH1OD
SGZ(e-?V.dFYN7BS9>I1FU;YG]VB??TbL31QJ=+cfId7,\PDVG+R^KZ_Wg4EMbK-
LY:.KcG=KZ9KRZ)AC6FY-;Sed1[SV;dWUX35Ua4BF<\)3ga-AGfP>O\T-)8^b@c]
UP#<(cN1VP<=bc2^bcU>K^E6aQc>GDDMVF6^WgeN\N_UWg9.OgE8IG=P>JXPP&V7
g2@(J0bSEQ7<V_@a#cF7K6?DFHW0&/faU<TW7EcSKS/ec2WD47af^eH-cAAT_]?Z
)<#>Z/g](R&\\ZH?]WHQf<B##[);[gUO,KO2/]I7SMSQ,[881R,]JY=cN)gfXD#&
T0MdDNcAT(8@EK^d4&Rf(P3O^7ZRMf?=;N+7=]=P^@Q&9=P@W7;\-TY1=3:D3ICZ
Z7>>,F-F]4P\=/LW;0(&9;d(a>D@e96OA2#T+2NP/PTM&F.<PF)<9^0B]<g1\8ZJ
+M7&)-^43/1;ABFd4CFcM\5Z)B@L[BcD->O>Xd^8_;_cNb&b.J:00M(>1KHFJC:C
8P3W&P359=Q(3KHYNXcR2.+\-(Y=]RBag1HBeM+A]DB\8,0HOR1&eMY9I@7#SMA.
NXX5J)b<:4G@>^7?\OBFKPQ1)D74OF7=1]IUOO:OFQFTf(573)Ge]XUGB,(A[,U;
]?-L(eX>8B7.1H:bW-4Gg8DKCLE0/gd<Xg,POcTFdW2?C&Zg^C[/F4GbV,NefP78
DPG7))bSe-T099FF1,gC5,?#/5>HW78X]I)?VF^e<cC6N.7^,,IYRCc/AYI<]GRg
,ZLKE=R47aWZE>?(T@VI2;2I8X)J2ZDUXKH?=9:G>U]^?\.);SLPOBIa:A4-(a3_
]M&6b>QZSR]TcfFY,-Qf&A0]HM?AB/[#D8f:NGZHeUbF/1Sga(LE^_3ODf1O]DZ^
g/(VDcg]=[RM1fQ=1QP2(2F&7\N4^+#5?b<c[4_N#PUIYXc1IL?6FD[[V2J#U;Sc
JMR;&Gd)7DR=SL2D<KI;@YM-RMbD@ZQUHMb./D(13N<@QTQ<FPJY\WL#&<NP46Z0
ef5c+c,E<,SZ9]Y3)3\XCJ_f=1-=UfIRfc:(R-g,#SJ1JTbfaDCAZbL1R8V(=04)
dB4=9KMa0OXSPUH@bc4K7&:T/J(Jbg]P/T8(-^/bM.[ZIM8IAN;W]RTP&b1D4Da3
520W4N:cF#b5aYR/ZRJHW/L4cL:3KYK>b79eC\\\e[K+Z4Se)adSJP,L@VEQ-S4S
b</BDU?L/ORHEGVOcDLE&G<[G<P2f0:0FZ.#I(EE02(Hf<1:Nbc_=8gE+T\/ZJL;
bCfHOLO:U3(BcWQB)C8^5fG+g-JJV8\ZN&SJKLUFNL;71)_#ZSb(/Efea.:#Dc]]
8A6f,>;XE<Na[3fA_AB9),T;?Z,7OBYUXdZAg?.EF8&Zc4?aNRfQM.R1/)8@O,SN
32HCAX/X#ZAKaSRO@NKNJV3CA/K^cKYXB9c64EQT5X-)>^PdeHQ:L7/fN(JKVgZg
.]?+06H.99;P::b.O7(7I4T[BAVB:XWQJ[5)R5<B_bGULF8dJTK13=LdBWK#TN5<
=V&;/b,_WGSa,/RdJ8Re3;ZXb4WJC=5[W6K_9ZKd&T8Q,)E@8;e_b/MU)ffQ8SS@
H(+=L_B/:DJC3R(=>^..,)WPfC<0NgF56>RJIPD8&PR2B;G&\cLY;=\FRWS157K(
]+fMW]=G>6dYMSO;FE7c@AX6F6>_7^a)?+#S0;8/;Bf_)fL6c82L-&JX17S\\=/Z
<fBAPY5;R_3&P,EUX+Ya>:P_\8A2_EY1.FKBL2+HILE)gTOgV1TFQ9U8D>:41ea_
+6eGXNH@CPF=X1bdL#F#Y9\2QM+ZDdLP2A+H(PNaP,=Pd.ZE-SR7.#)&ZR(_+g5P
R^XM9e@E?T6N(\3.HDS9:_T,,HVLTONU^I9))9&F=-YFF-FUY=Y.dLZR)]OH@&_F
8;C_5\a4CPZPaDPBWI>AO#F3477/->F0+OS37^_1FBbS2fMETcDQJYLQNOXQB+^G
M+I;fL>c0)M\@SZ9:.?OE#CV&9OC5#eIE_@a^JM+,/LY7<LKF]/AA+]\XBfA/5]/
[VeCVB35)(e)3I2YWN7J_]\7M6=:V&K[d6TBV-/)cGOOXEHTLR0CMPJEPJBG5d3E
ScPb6O<A5/ggVYeE6N\eIDCDa7+2XNF?,]M4cH9GeDcCD34cN:;bcUF7V>QRW<WB
N\/2,LB5=.6<6T6K175<JD<_DX\#[E]a3B+WK<V6[0UR(4A7@fX4/YP9M6=/[\EN
X4E7K@]M.eU)+VSJ<DZEG:UC=\_I3F#U&+NL8FaIOY6E6U\936;U,_M+TfQK,g&O
-;YL>UX+KP?/.FK+[XfJfV<7M7QIaT#47bQHS0UFP9O+_###(GF:Q&3VKQ\@@5c?
3:Sac76@[(]Hb+K:1Q>YW1^UFR_&(.cP&GSId#ZZZLG#]AH);6FC3MW286Z3Hg;V
7J<f38GTAFAZJ0R<RUaY:c#<XgWU9+M>M_P2X2552FF>,\THAWAHY6BF-aW9HT.Z
;Y/5VNd_&B-U/0<91\a6+[O_69?K^Ig9;S81N^;FW-:;=,R.QU^cL+C\\D@&,QgM
>ZdE[W7U(fc=Y5dG])R.@3_/&21H@[]/=b<>T8d(NK8&dab^U6+R5\S+0O8(V.D>
=d/D@g,/T\OWQ#RUS\3bDJ/X0g<M;5&HZ0JK)aY7.<^G(.7=_L6[bb;=dW_NKYf;
a6S655KOL8R.X0IcPT_\F]M2G)AFT8VVf[J^b)DK+BM?==de8D56UgSXH2UAC(\G
FY95\P:S1ZQg?_5)1bW)B9KTK9::0c4A8@Q-OV-Y&P:T..XV7W9MG)AW3FP0P66Q
_f+U1Fa^Af9c_O,PfWM=/V@?;QMA862OEN1ed(H>)9EU.SSD71QdM<gg6,B>V_)W
W53DMGBQ+2+aKA,2Be7,:HL)W_/ADaSH_I71dO9Vb[0HXH_SeI7,H=697EC=#bII
].H,YWgfT_A4XD:2UMZ?I\ZcS0beU?YaPf<3T\2TAW-BHL^a:6I<agGH<74eYW0E
=P_BE0e2N0V@)HHQ6>0;@cI_cCc20GOQ=G^.cA)(EVLCOV>WFK=/-LSH.OWH)>4@
;G>Q^=@b2J4dB7Z?&#:fOO&0AFVFe\\(8KJ7g(gE8Me04H5Fad3d=JDO4KE^@/6@
H5E<.U7X@^c-dde0DU,K?b]VRQG:a;]/7BR<fQ&^X23VLM#UBI>g4F=WF;88Sb[C
c+bgF-<c88N^/NQP1]OB1T3SN-B<7P<200C6-8WcR.[<PEMa]e#F9&U2T>OI<,>-
#=#AM9CeKVCXEPgTM>gC&=O^?6Qb.U-UUO1^F(34V<NDRMYX\/0bVPICaNLA32(6
d+OJK;A;]3Cca_a&Bg>;H-bL&;4eL25]&g2,LM82UD)8G97O7RBcGSb-a^^IRa=R
T,S_#)(VVD^/cD884,aCT25M50S?F22O#cW99cR6HQCTBX,6HBWUOQ/0f[dYTC=7
NdT919Z^/>8Uc#_bS6B]V)@O\;_g>7c_>cJG^YXb6;dDBH<P:->G\RDe4SaI5e-e
eF-.2Q/NT>13(5NQfH<TR[[Sd1;<cb>4P@AG7X558H<M?2,J#:d>+?g_\^gbF1X&
+Q^e&XZT2<4F_:<//&Y?#FY4_dg>Y1L?-)(e/I(daX_MIN,Xg.;L3;(<c/Z30W(1
V,5P(O<HaLTS23-g.5Ifb(5Kf?>T;V\-&H6e(#SH/J(\9&Tb@V7Y,Z_a1\:Z9f+U
8:+/K[M9>3;4:9A2I:3?\3GVM(64KaSPTO:8[O0@g)B]03/cRX#e@dPg/5:-Q2K+
RURZc/XTMK&_HG\@^I<^S[?]AZ;^]_WKBJB2c5d@=TIdMd;)&B?.9V;HQV@/]d^R
6[I-))+Y@.3WaH-7Lb(f0FCTY)35C@B.4DH;)]X3@F1>ZCSWSa\4:Ub-MEOE3+)F
G->_.1,?ZF)7PVFO=c:LD7.Lg9R>,,J6gZ,>TB3B395?P76/\_FLGY/N\\Z/Ye;,
T4TIHL2U05XA5,B#\C:U=.f6eTc6>><0Fa22E]WV@=]dGd-)#9E,8dQJ8-?(.(8e
5>[:==UBg1]C,KW=eR2I;c?MfeAO]eXdg^.?B=[V0JJDL/3d]SMK:9.U.#2V>MMF
[f&N&,C<=[8bO3OF<LE_Ta(7E0\8=XX9[=J#c70N>(;g4IMGX5)\-T:748dCW+-d
5YFa>cb^RDP9/??(B4eTaabSBA#aKU9A(E&=F\;_>(2VE^G7-MSI/g[/PF?P7d)Z
H#4(ZXV6\-5KR)@DZ<B/P<9CHM@JbA#T-Ua0PG592/B>:>50YIe]5FeXGF^G_7)X
#+Y^0T]baA1fXd<AX[c:321>S&3=g6VSEN&5NII<,IaRP^C.=KX(O#c5;R&-M&89
W4fbM]TAO>?:0?d3A0NM\J^)9e>MF>UV1R?bAbNbgMHKWIFP2)W8HYR;dS(7]V(G
EM06:18A#M-+Sd_,d0VB>6ec[F)fc..Q?G47PI>HGT_(SJaa=dQ<^/&(^dS&\N(4
/J?Z<=E?T;?50(TOe:&XTR720:>f5bF)W8IQ07M[;+9NAEf@4C;K^71[c\?6C1_F
.PV1(5);>/PKWe5E]EH1I?5]QZI#VQfJJb/2ZM:ZYdC(VZZT\g]#];FG9N>GIRB?
aSOL(U[_-USg.H:RG9SQe\:8fACa9NbXDf?INH-<L=LST3\LU<X,1a6b3_C<@ASU
M(G;^37,W+d8<LLPM/QVS.@4T1N]7F3RW_d^>aJOOXSZ\-SN5(a;CI+S)0T32\EP
4b)1H[LO9.IUW:ZA1V3GDJNCJ3SBD4]Xb<VDZe]dO_]-d)e8H.2/V?F,LIAAFTM]
&KdN^M?M6.=Y5C-#>NE,a:A<^<^PGQ,TPfL21AO5F?9]5SRXDe]8,C,:Y2.T0,eZ
(51(MWZWN3?6832<Q]?/X#WQ9+RP04DBLJ7RU?0Q.S@e2U?U;e/>IL@I.ELdbE4d
F;GgT2b=EK^JbD5?-CDD?NXKU@:K3e.)U=>,X4#W0H^O3#WFG\eW@Tcc3DW5_<BD
\9)XCGg/\R)Y7CLHeW2#e9#DL1daS;>b0V#+^G-aIC:eI,0_WI)V0OCO@MQYP:DV
\8bfUS(aLKKQ#e>?_:A?F=@,Ab/YF:BfC]4)e+JfO&L8TXZHDda+^;=X92\2MRC9
^1MA27&L]cHX^YVa^YTB.A1IcPYP6R>&2HVg@,Z,_A[^eM<)(0WcVdO0.gAR:/YJ
L?N/X1cg0/5SY1[UbA1TTS)-c]OL2Y+-H])UU\W]X3NIeW\>70(#bUP2FNXJdJ68
F:.gL61PQ\T0<@f.&7V0.aP3;OYJVM33[91?T5DZ,E2gdXWb^bdJ3J/\#_D56,e7
7MNM.>O6H4^?D+7a6C2UAe5;.FJ_2(^Y9^d](.]9?=[MR&?90Tb3+W]&QJM8+<96
3dH+3C3K9L)C9<+.F##@IddD;663AV;XTF@b^#Y,QcT]VO;3:7JMYJ@-J/_.aa=:
#3M6BC0J\A:?26,>(YHEU)/W85)K@fC=RgCW6>fLb_H6X#HOE8\OLVCF83MN[&T#
2^O>0[aa>&RL>gX/?^g,NP,OX:=GJ3]BKBa1P(V=ZJ(]gTPECV?D,Mb3EFXYT:4b
(c?IBJSg5-V>De<&ARVNU,dVQ1adJ:OBFYVH_?PI:SbX4FeSKKLE_4MbO]+B&^F9
.+>,NLXOG.Y4B3FTDG(:\=\NZ4/MPR^=P8ZDb<[^<FDR48&L47.-)#Y#(]4^,-]T
X]CbQVVR)M.9g[1Ee@1(F22cPTX5FU\fWLJ__O^C_OK.1MTR?^/0:OJEV&#K2d66
]GfURSZL@&Z8e9FaRLgYSa<IQVeDD3L)J(\Q+G[<L&#<M<8D,RgD#.WR[YIX_Kb=
H9J;]AP8NQW]ZT;M1D-X;Xc9<Y(fgE=3G-E?K1D68@.4Y9HJabWRf^>BM7;1^Fd?
DcH3B)XG,>H7TK@&WYF6&Q:f)^GUYAb_,J3eB;ec^SP4Wa,AK6#,]ZTOY-e3c-#K
4+84Tf[Z_J?Q<(GA^aE86&KPA?Re^J91#,]9_,Z1W)\H_KbJ;,<9RT2e6.[+Wf7L
HR.>]F&YP.\9Pb\3XQJTGNS;X#XL6J_IT.OT^d^)cP?gE:aF#QXFD?=(6Q.<_@_H
GWAEAQ6G:Ua@QD&2-gbNfL+/#1H:a<18Na=Z[:f,\R\bb(.CMLfE@7:#1SOMd@e(
Q#MPDC_+RD:;#IV;T,&U^]A1dCKa-XP_INdba@4KUF>LSQc;_#-gMNZ46+\[E-B4
)+ga?V29fCS_X?MF2K^12bA5:P_QFDP=a>d/^@cP)a<1ON#LLTe;b2@@&(C-?N?;
/,Q+J>e]P.Q>S;?^=ADBc?LQ#bKa^4aXH,+_Bc1@:>U1RD8I&1AI&@9\/NBP@d#D
F1gF0g-?3+58-:ZNRT_(>\a@Ka4^Q\f<8^I\e1_QaR->:6:X4JAU@Q--a2[V#O?F
6aUT2HJG(4)/Q>8BJe[Q,4JJRb:0-=]:DQT@Yg6&S);QRS6XDDEVD(agbWga;TL/
PFde;2BGN1ZfDMd9e9VQTXf0#52Z[H/4-O-ORY^K?8g.?Ya=C^8B+LNM3M0UQ3\V
FF/?6_;03B#<8Ee60GY<VAGXI12\RJ;gRO;?bGIF@_NDOXT-&QNK4@);;?b?2W\&
A([T;Y1S(<LYZZCH;C\gaZ9MF+UTaB>Vf]aT))225UT>8a?(Yc#e#XU4=#1]TZ=Q
K7If3)-0WeOVgG+;<MY=(5=87LbL=[3V?F.<@@aBfO/H;8RJLP.U_g/_-_fdBG^Q
C]#5Hc5d5TLT+FG;_C>,9M.)V52#E,gVPF2>b0fM5]7TcODdVce1_+gHG6[b\^MS
b?e5-LAg_eAQOb[EM@V_cOM<RP3^BELa/dOEETdYT>_Q:U1e0EIHQIIW3.Hc=6:O
R/4LJ>MO9S&M/Q;BY^D;7Q>3/@<=]\IA)H]88F&R\7U@A._4+eeHRTO(dZ09;P^Q
L[FCA<B3^R\4+I9Pe/fJ1SK_;>LJTe2RfWOfF4.+-D@-bf=]A>K?EJIa;aS40R2_
_MH\gZD@PVefY&He3C#fDa0Pd:2#F83N=SR/-4I3>b+Q]Y7a4K5UDO\>N-\F<62<
FIEE?aGP(-SaISLgB(2XDWPV@0EZVN3VP\-,D5gQVS:MCLe.K+:,DTeET9WE4f+;
cE#4c-H5&S=?]_<N/Q_7+I#H,:0&Xa85IZLC+S2=eYf/;-Zd_IB6,+HFeLL;+<Xa
Ag#a3SC,Y,)H5+VTd^R>)\?=7&7U1T]]RVMD8LR9b\5HA.P(_YER]EN?JV2/)P?G
H;36?f.+,GcPa8b+EMe5=N>]U4YG4]O,8P>,]WKYD1@0?BEM7:^C>84<-=@d8f0H
e])GLUSL:-=6b;PEb&R5X0g9K1F8&,2)QQab3P[3]_/Z?(-DgWbW+:--M)),1++F
DfC8GcJd.YaOcNUDOF\W[L4W4<H;-\:#d24-H7<4/@Y\P>POF7C>aL@.O20=@/]]
R632320Ue@/)K8-&G,7@2)N6;(T:Y7V:Q.389e[(_SXZO(Y([V]85cL&)XY(WL(K
,]&=),(S_Q4_bR.[Y55D/]PVNX&5<JQeH^><6_b2&_LH>[d6\GBNdK.\gMW3VGA\
@L0AK0_MPHSc;#\NVKEbb^U^_Oc\4HY:NMAKW;ZI-LG1NP[0Z-^G59G50>&86XXE
,#7U[=ca_CZf/)[>VL3bAdDTZ?IgbT/>>=F?d9-)?;LPE)F,2@eX:&:)[Fe-:\gH
,]SPWR)KCA2]_<&@]P#N]L&cV1FO80FaPB]CBCS^K5W9T(7FF]KVEW:=8],&VJMN
6,g>FA<dN#?AF3XZc/@eXb81J63H]A)L4]TUR:20D&R371;aQHd1X&@gO;KJc]bZ
)P8=CXW7=.H?[Q/1@J4DP&3&^8\L#)SG.F/D4cH[3[;00M47ObZW(Q6?F_c/:^)D
48B#Ha,P6.&e1?MT_/<K\&^N,+:@2LEJCc,b80<@NecD/G=?.N\?9[,W\aeT7QRa
@#BgMJBE0FTK08XK05L1TR?A;8(ZAWCC7;BKGcTAd<6T[8GEQ/JAY9RC\[V8S.cd
^3]QE,TF_A\QEL]UM.W0J\ad37Ae5S/8=9/&.Cb#c-O,@5]Jff:+<IJ:FRW6_c)F
44I[;&1@8P@3^LbLc&Y;)7.=.Lf7Oe-Eac1e>LFMd2IZ>AQ;e?3B^6-6L6^YOKe2
PL#Vc)-W2&0da=M-e4[T;aI>84/(G:@H(4?=cR8E=f9a>2g3?^dV[9]65c7gKQ=D
;U.Z-94?RR&>2K4+JgXCCQ\Ma^:O#2AW]Jb_F?RM(;eMeI7X=H+K_5_UDeC9B^_H
[/-c(5H0-E#05).IO1Qe[&#JRG13BUPQ@OOV]<1dBLC76-T1Y@?a@Mg#-E]9EK1N
&;2:]PJ@I1?N?caRXNDTcJ.=3/-eH7YSgN7L/^CVGSZPMX)Pe89D>DG(50&1OM2=
N3d8BP^eRO9-OUR:fabQ[+L<ceY+C,4E=\M]M,bd,5;-^/J:),K_0eYQB6Xg9VF6
T4BW>003R9dR&@;)>1_JNV1G2];039>CXX?XWQ_5D-[1#>G>#:5?ZZ+BO^8=4c1A
#58P6:F_[2-9)9)eFU4]\C&CA>VJ(e(@N85a#HeB^&PJd4R,B)->P6If@V8+8\=g
T4JI.d;IR4RI82VDUC:/783W[e[JX_?_.VfSR0F6Z<DL81YP74&R16_WH5Q;#dA4
&C+F0:BODTCKB8eJ)/\5FQZW75^.=P9KUPI?6.]^Y(eCI._9@g[;c6ScfS(\[ELC
\V@(6F28KGN\)4.OE,5(W0^.3>C^0fB:B,QOO;.W6(F;Z]TXIF^[b<H8\LX(WXD7
1CIO]KOAIf@I^1_G):ae\_3.L:;AbfEeW4J.M(@],7JBI]dO=)\<STZ(0+5WDM1c
TDNM)d?(;_<<.eCW8QPZc\:^d.0ZfOSR^XgWF.f.0+/ObdeOVA>H9H9?V]&X6(dN
e8Wg@#gK1<(=_GdK)7cgPC-/6NAD^b-VX\IJR[dUE9=g3,&PS79M_TO.IaX(=db;
Z.G^(4f1^1ee_VKe.<)-X)@bV@S+NHOTeSC(U+Y3_PHI<1OD9<<;SWf5&NT7L<:T
J)1WX)U2d61HbZVRJa=U(T0I;e=EFY6KR@P;CR)-KCL;+e]Z2Df2\<.1WTP??9;a
G\?IWTYC-7&bBENU/g3PafY(<9LE]V=A58GJ?XdE<XSBbIBSc3XQZZ42=SI+e;FO
DL>F9AT+=^3<3Rg@BcG59b0dQG3L40__(]]VMC.V3Nb]Q\_ZE3D2g^]MHg8cKdfU
0f:eJ5_6Uf7LG)Q.9_R>TJ>,Q.8JQPHQPc4RbH:\eARRS7b_HGS1O^O;0a:WU1Q?
5+[>GD;(-[a4PSC,QX[W(Gg2LW]g8D)VJ-aC+I>(AH8aL8#I/&b)#H1\:-^+XW4N
@8Yab.-V?8\,B:9&XHNTN453P2(RGE]gDg8,Q)eWP@g@\#&=2;MODe#WPU3E9;]I
2C_6#d_M8WD4.W7:daa2RUS5:4N?Y1&SV#gR+##E#[O6e;9W[XDVKEFA=,;)gZ5P
TCPe+MR0PDa6#fJYBR)2:^?#_eDVEP7FER<W3eQSW/Mc@^35MN3YAZD.@cg;,@#?
&Sd+,3;/.C[^GWb6Ze-FX])JPJYe)]bEBNR?b4;;dBD8PI.8gAO<cc_W=@;1W3-1
.BX#2gSA]ZAGB,(G=8Q\]c9:[08N/FO-c22)8-YNR)ZA<aIH(c\.>(A5ZD9M&91S
&R5[H6D4T\CP546BGA_?aG0Ag/L2054d-6?>N&O]HYEU15E6;TXOZ+]D^BD/QbM1
H,P9OWPVO.9D+0(].&9CI5KS-gBKU1Da5bP@E_IaZDaO;eMV:9#<8Ka/P_R.2Z/W
4G)8528QL-TDS/-e5].a:g6(]@<2FH=Af3O8DZ_fdf,0c@(58[N;b3:)4f^#:)(>
:O500V9C_UZ2<Mb;HRY?_(Q&b^X(07I09]\,Ae[0G)5a,O[#5-[c1--&d\EX::V_
PNIA7MBV1=J>HZd(cV6MZEW>+5J[4^03C(f^,9&d?:)82)0dO+7>R^6[NIcRe^\8
BZ;N4[=g<R-[Q=DS;H.TT[B]N@QU@OIK::G2KFc;ZKKDXXOg]Y4BA3PH/(HQfCMW
8>5@B2?<g+Xe;6OR=9eb=80CASR^SI.fX+0@11cgbHRA:OL4QR-=Wa)QJ)S8>Yc&
G-<4=cI1b/9AZ[@02U#H5:<5c-XNIUXZE=Ia7(:7(-W>A:.RVV(YP6KJB[Q57=LJ
1_E^#QCfGWG([4[8#OM4:A48:ID&YUJ+NHe&YD)ULCXL@@Yc4E?]U1C4R1:,f:Y4
->6\9Z=_DV97M1Wb=HM6?Q36#E/ILWD3:8IL3)RT052LgCg09M1(E;PG74,0f#GU
W\?I1Z/OSg.A=H.F0_-4JO4dAMK\0AA.+X1V9A5M(MP1U1QV1cJg/117;?^;ZT.g
FV\F<cZf-=@)LJBb@(4DN>&WRC5]P:X>@27P9g9I[Y@[O_3,,Pg+8b6EEY7DXcIV
CSfF0\Y2a5VVL/PPUeF>HP>R;D[T>a[?bLVEWgFP_4\0;aQ)GCGJQ.MOR(01E8-=
SH79SBLL.,6cKOFT?3XQG8Y[IcZ3g\2@bN8PXcGB+4#C0;;Q)(K?>^bR@[LTaaKX
KV/.O)9.+^6YIPVBT;f.eHTZW._(6e&03P+P.BR#.U@PE\8TNK#A>+TR\3A+94&2
cRW-c)9JO2DI84)SVC2Y(KNWQ:Z<2CZ0-5F84@bG?>BY1fJg08&)XI/7E&N:EbH>
<7ZR0aY,O?U,2M/:c_?P;?=2<_+JUSF3@b1eIBGCQM4<3/ST54V=&[0ge2?6,.c\
@AADcL)ZODEd0/&D)U\3LaD0N@?.5YA+8Q8Q:f^:.IY1X/<?<eZD)cA:TN\MZG^(
/(c</b\KO?^VZ_9AX0W4#;&\A(\Saf3T=LC6E<XIf[#QMY<XBB?9(GS)Q[D-58/@
;&N2FCDBS1F5(V=53&TB&Y8(H.49S\3;\0bC+4O11X?X7d.N<:_TbQBb,D_G[B)H
=?U?GC3d6>E\._JD=MK9..03d_@Oa(O1HB/c:64RC7Cab=:ALH,D5MaL@>0Z+Y^B
P;dBOG,>eU:eN;R^E\3\I,I29Y9VUH;IHJ,P76TW1S5V58ffQKADeR_:,cP_ecS2
RVQP.AP+)T&If+Y7)?9+cg6Ff,,@KS?e7_]BdK;0RAH/\ZgD,>[NARZPdgWC2Uc9
[gg=Z6bDY#dQ2#&Eg8UH_aMg[4<AD5_@)[=[H06(M(PW=AYPA^?gY4IM?6a_05(B
-UAe@\AUf2deYN&J2@VH5D)N;MP8QXI?@_SOB95XSb](#^5f@G7840-GOU2_DL<P
+c>dZZGBXB6ePVZ:fd1WNNYS_32M(CPDd=N5.f6#dM7J92CVB@>cdAc(&a^)V^[E
M:=BfB_2V_-W7FP=J_<(K>-OF?G,TeF&CGTM5NQEG[MIHUUR7LMg=8ZCR3_ZcCHb
EfJ4T7PUeY7c<T6H#fI;=ONe\g>4_9;?=<X9_)OL<7G^&DNGG[2?1W18agHIbS/.
YXL&a/7=I&EPad2E<KD8&(W6B[^^ECH.5Qc88EY<e(_=CbTQ9+9L?8X<(LFRaLC5
Xd^Y;ZUQg(DP../-])f>(MS.UXX]f0,,DNEK]W;96CEUO]D/dQ<XZ)g0V-BA]abD
:E=?_M,d1\+UWALV,JCUU2P6HBE?3V?FeRT?-1Xa\(XHfIbba,.W=W_T;aZCL_@B
H,c]49QF?7J5=P+KCg^.)cFL,S0A+>A->@P@31GUWXPE7fZ^U1X03a1<QY,C8bG:
1[4SLB-#@Z#B/4/cgW=.6+\P\^C_0I^@afb[cDV+=/5ZLLGg#,g//./KeK>#<aE/
.abG(c45;N&3(YLHPE+3&BbV>+O+#G^9)ZEQZ=>E_?67N^g.a+T;4>U@-ZC5.<d(
aRCAHa3F7@^IF2K0?f;#g4,#.WLNOU2M=2+6-XTc9ZT9DD=\EN0]#9I&V)gTT94X
H?MO5bDCDF=IHa:^M^)NJBQX&e4?6@9?+.=ZCB#]P^eNJ.:.gBR()5Bf2CI6ePHL
8PX\#W>WW):3+?gD2_:Gag8HYP\<1]-cE^dF.Z-(@SMf1c\K31KH_[T45?>6FNa)
:,1D5e?&C<EIK97KX@(&NB1OQd^G30V4MNd=P=eEY<d(.>T]/[\563/UHJED=;SZ
EcG?:]F9HTJ+N(@c73JBHEcEg=M66.gd5,L)I@;<#6ZDfFM(<PW6XgKQFdO#V6f3
J5L8^A-61./(6]76.G>]0fWRPgR=HgdB1G@aCI29FT.)958fVV;#Mb<&(56V<g7=
7WZSTUM)&7Zd6S1cFUcJ@Va1X?3W<2IPC:;)4If>Y2TH5GB286C4S+BM_4f?6>54
^K3<HF,3MFfVQ[DFWF/]>:K_BC\#F2d4D9^Q0=c9bLcg\P=FDZ@bGCd;PTe#c/UT
\9,/6DWfC?^M\R3DQUT#;8GgD;[M8WdNPI9#054d)4,Y>>.8EV(>.X)FVI(V?WDK
(2B6YL5^:W?TNC@c#[C3(4e@^baf(K@N/Q71EM1RIOC+ASAGP_UL4IZO[Tg;6cDc
H@YI?I2KFQ\>&Z:T[a,WD=bRIWYXI,c@)0J[NKQD>&OR7BO.+c:bZb@,EOSQf1P[
^^Wg4R9N_dEGZT?Qdf+;MCX#]LS&YcK-D#X#7W&b51D0HaC0/aCWMKYfM]6AYWCX
OFHLSf&Y=B.(O+(>FEF^GcC]AbOf2.=d[^/YD50=dH-S.^O0Y&;ISHOcG4GL)8@L
fCbX4:[..D<AYL64(5.Y4HgJ5(LEG-#:#COA)W8dH?\5C74A,9&0fIbc_.dMQabO
K:W_49/R+[\\8PDKY1>#?P_;+[=O(,_5I;OAbI5T]Q8N4ZT3Z,Ngg).V[<C,RUMV
1#BF28&a_UF>H/=P2>f3;bF#SV=g(dU&P8HScU8E=>&I,M]EVLg]XfDR@^BY/3\.
L-f9WD>a2L#Q@dQ&,?TO8/31g,72Z@.5BbdOIYOK=>eIK@YSgH]5+5A&\:?RT<R8
ZcR(g>I2E+9A=4O&9:^f_RLYK1a6JQ+V@XY<_B(<34X-EC0-H7YCZ7_W6a]E3H.B
&@.<M/Z65>Y,X=JS-]EH:.KUQKF)+C@\#[52A=&XN[]H2&[>>e5ZGg6W+.AR9;YV
1aZfA#,KU2aPHfB/41(E9Y81FbBF<=F[2+SWR7Y^9BVS)9.TR6F:Z.fN+P@F2=c8
-C<RX6;SQ^[LV6:?VLHKW-22?V(L6a/XG,.5]]U=]S-?7E6=?F6]FJ_.cd7bdQ,(
0(=5,\H)Hg0cWVWcHOYHe>KPQ\9:.dKL4R0[VN&PNd+I1U)[XOYH:P,D7MYgRa&=
H?DIc/4<ABd_7d+?TBJ?-55#O>0LLb8^88WgWZd#@;D+^53^>^3GA^f5:8bHe.;c
gU_]2D_)S>HZ^IRd8a4W,J/+)KWa6DYeZ9L-T(MH=e,ZaaG7QLOXfI.e&2g+P&g6
FD&.#XD&3fE@V3P&GS8X5+1e?\O\TY^d49[-PE6N\^;#ea^K=HaDeLLFX@D?V(JI
dH.X?MeI#-e_bU7EH3I3E4SE4M1&NZ?9/;F\KS1I#S;-5P9]Cc=WQY1HE7ZMSb-X
Z<&a^>STPS\&9U,)4\[6;)G3G@G^Ee.70[LBBd)bDY^NEe1G]TTKC[M<2&P>KNg1
bHI,4@EADEX4XLX0H=(D)8C=0??e0^.8A8[,JB\UZ(UQ:@eP@XF-cH?0fgYc4>7(
=IL&WE#SXYS1-K]\9J?YcGL\GPS:e?;OX&b#/gP,f+Y:HT1ED.\W#_K?-1\K4FEM
8E<;BH7>F#P^XKO.T@2ITICH;X:<c7@DQCUFDELE(770I=/)d(C@Ee6G2A(H,9bX
]TPR=+V[Bd,6[H3TB0HX3?N<H]e74RIIO+S7bIJLU-aQgROPQZ&[HD3HJTEAAF0A
4_=RKDIcQLIBbD#->G.#PL=:J(,ZDN]6fJ^1f^76&K]73NCQGLDD76EQc.VBN-BA
?WbYCIIF<e/5#ZQHaXW.QGgSN##gT2)?C1Z3Fc[:11H4WCDG[V/LcO#>e]KW6bVY
PPN3ObDe[CG[,PR;]2.60\eOAXB9+TY\Udc@T/;J;]+/,K2e:Y7fHb,0_N:#P^5P
X9CGM2L=cZU?HT8W3Ug];a.#M=S]4T4&VOLA<]K,CH?DcUVYG6+=FDgT&UDY27#X
:-J)U?b\&)[OHUTO@.V,/5SQ/?XdaC1]4PNW-042+R6ZGG79]W+6-Tg1GPbX7VY@
##\T@aD&9;D0e_&\bafR2?[@<?RH2(^3REf1T5dUS#_@XaW+R:]#CP+B+0e(5F6.
[Z2^N]T=HK8K0+dbHdP;20gZfYG)f)^8O#WRTQ?HW0^;eD9K\OT_La3@\9E(>@@>
-F:14gP]C-ZQ7+gL.VD(5??3;)0(?MT\4J/2,^.b?<:,1U4A/N37HdFgMf,IU9SH
(XG,..1Y&XfG6_BU&MF_gC]-1<@c;Z,IN+.YU)][/7UZ9Sf:X@[D(MfC-IF.;&&0
FPXL;=\X50Eg]F&@;_d0)aPgeFM0J(A&\G^5g,QD.AADV0dZ1YVW]<B)PN<.\c11
3]U9C/&O<ZVPML/X3XX1R,T1<;<0PP)=FNFC0R(aE:SIH&e1CCKFVIdaPQ0XG+57
Mf2)VZP&\C?X1,g1D<O-0AHIL(ZKU#K(L;<QKea)AZc0HS>E(9T;IN&]<_e.c=Te
7?AbgLT7e+OS+.^W3NV7)Z>TJM<PHNT9VPYCc_Z)MXZ?Oe@gGEd)H(FEN/G6Z)W3
./:B6C]4J(=TB\K-@P[U7L@4;_GC@f;P<Y_=c.<:G8:?6OFFPXAP43C@Q2^#ce?-
M0XRXc,Q2gf2,^IYaQW]:#PPJ2>LQ_<WRW7PdaW#0>45N23+06E6^#<5U6?bRA]Q
aY,=;(PP5?VdDC/M<H7M.P0GM0N,4[<@6/?g1YN\(g_=G<Q)c?)JP,U38b:/HALe
6S40>fARYMJ+g,X@UeM62-P>@Z++#?;I71MKTU>P+HfW=aO?:K3.]#9TD;<PZc5O
]F=M]86:>NKR)2:2MR1((gN9>HC+,T&<<I8A@WLO(Y>:).=;ZKDD[N>,Nc<U+g]A
B@96X^N]FE7d?7bf&[Qd@=/;Y/9B2aPZQ82IN_1^XJX3:6@Gc,2.[3ec7FV]6+#&
fXUc,E9JZ7=6,\UEZPP8L+(d#c4#WCHL7=I50.71dMIA-Y9C[=Bc.OgEW4KR]RB[
4DbS>aOUg.2N/-6PTDFY[<1KHZYJ\Sc^YPdLA5LAPIM2@)2IX)[)Uf/5JGZ7Ha,W
f0a<#>7g#PceH_7@5]W[L>dH@.G2EJ&/9^2DW7?MKR_Jd^AB#CAU/D+Y.J:SDMB4
6fOFPHL#5/?;6]2.=DXS29HA7RKOAWN]6#6X+fAZ[<\L6L_[d+U&S6Ifg7O@-Y#+
Sg+U=I\HaaBgc731_-aKBE([=U5YMV1C9<b33?56]&FMLOLdI-)Q3VgNW<eT2;5d
T>I0Y^H1[@DeHM<=@7U2@_L<W:.66ZN_LK)?[_>RLIgcFFG45&^LA:SUX-,+DaM5
[V4^ZS)=C;Q\7c5\+/2B&#ee?80HcX&8^)+2S&D=PU(_L.>7DE[LWB^7R.Z>GXDU
#?+(TF.d=,Z?KL4PMgGgZHcD=BXa_GNY7;(VQ)4&a+aKK850D0CK\?<)+1Z6UAg^
KF6T:><P>>+^bOR[0XY(51<,<[DO0,BdYa_cHP.)V10?2.VD4eXbc<(dV8gPb.M]
.fM?=CSH+[b<3-4_#2]+24?HS42_&3:cM<::8LQ[5cS@cf?:9?IJ7J\^D5&=M7.]
^N6TTQ>_NWHAFD2[)>c3-F/VSG,CS(1VOc]8C92Z8-O1JI0D:1V_68H[=CRFEbW9
VZf?Z@3HeMcVM_YHSH>c(&Eg<7Y>>B5(ZFAQ4NG0Q]I/6:X0BdULA(&O9-I<#TF3
48P6;;A75NVeBGHVOR-7e\F5LQW,V<Hd>6fQgd1#deKA]3XWKg6FP-T-&Q_,_>R9
Ea60:J[6JE8PQU(G/R<8:L].LVU.JX11/=>7;7W43&_:F)#&M[7Y(-g&WHU7^:Sb
DTGJCFKC5D.4O>A2M]_I6]C6d1)Q.a0&K),@/IC=2P15IN&>:gFB&._QY(UM)=0<
IgZPC#V_;C:</9OO4)QY6>1F@JYR>?+g4f4);Y0eX_+9>XbJVEH&1M5A2QRg9CXR
WO1X^S1)U:fGUV[E?XF[a:f8D^OJ9>B8BGWEHgNQ,85X/ZML2@A(YW<SK2+(QZ4+
5e8e2:Zf=5M2,a0>#K8V)Z[4OJ+^4M;&_E,N#-T?><#6aD?YFAJ>GDH?R_=K5X1E
VW-=8#?&fBB3A&dHFe>/>O&e2SN4UG5(cNcNg+)5?3PMdEM\A_b7^=;]=/U+T].@
@W96>C;2J)\E\,,Fe^^1ZB>SLKZ<W+4)CdSXcBC<f)GKDUZ8PPdFKcCd_6J_8;_/
1DFM1SPA50636U:Z=?Rfd<GRVG:&gYKV&UMOgU[,PE\U[<XeR;F9NHfWf4=f,_GE
+=g60eTCMG?Z(Hcdg;ZdK[I=cUR83HU28IGNMPP,Dea5^gBQ[&-6FKa)H(P70<IY
+<-Y1ORB;f=E9dT]c^>NCN,FCZIO7R,<2=VX.^f85GAfg>7E[WUcXD(V::(,J-=M
+5]^896.edO0F9<Tc<(K4NB6I2,K#^3CVB.,8a^c>4]eS<edIN@V8L<dWCEd4b3&
dNRAa0afCTUDL&e:_H58-<F#_Qc1gS7BC1]^cTZ-&YNQfg4C.RBNP47Y28BN=03#
M3L-I0+0bU&a1b36P6FVLXGa/NB&)?RT)+10U_[<4QT@Cd>9;Q-IUQ&^NabaSA[K
3C4\4:9.b+R<GLA.OSC8c5Bf9=^(L&OK)&NUPbW1PG;J6]BR.,;9T:GFL@B^J=<g
2FCg+eTI_P8[Q9(UN(/_:]TC).BAA@c63^APdfY:GVdFe)LODZAK<b^JDfeYBb6f
U+dgT5c@A_,A9A)(^cUM,?T7:,.6&W+#B2F<FJ&D4Y-g^\M@-YNZMJ),9c-GXF5Q
I.RS<.CaEMJbM7f/E?c[+g7S7HB1(LI3>)/^(7XC>L1JH;4^8&PQB8\3.RFScbLc
/SRM1^aJR[#,)UdNZE((,Zc#LMX&WcU,MS4DaMe?DKMV=NOF:EW+W4R<,5a_SU?-
GGaGObBgWQB:]8:g-]CQB/05dH7D>abSCD?M;9^?<X-3S48_0Zd:FYJcNPU)bI04
,K:D>#-a^#QfB:BIT.45[:)3)c<Fe^d=EU33J17J5F?,69J)U6Q#XG7eLA84)D;4
1-)40]>beI0955SRIT3&A,AI?)^+e-(>J(7)dQM^Y4(6Q.Y?g9JR:6G5?H8PX).W
#7=gf(KC&Uf&@XC5)>+/.)U<Bd\^R=@A)X#RaE?XLd0#+FMS2SI[#Je)8,<#b>P4
]a0GQf,A3a#d2U/5AUHaI@XHKXXMOa7YfMRERV)8GQ:HbVNOJ\_O??@[add/I)5=
I@(6Bde#@cT=UA>5>50D>+^F8]N)N3a+V(]@aW>.HC<>1_>WTZ/HQD,SZ#=@B,Ic
+XG,>66b1T+:.S)17&Md->ME13S^4d1O\H9-63T>L#M^Ka&Z7T76WN)((VcV<8(;
fcJXZa2<f1&25?(6;KJQU\)(\8P>?[2<.d8#d0GL:-FYUFWA)<d]V528g>IASOBd
#NQc^G\90fFH58&XE?\98.1UFP]XX=e>G#=e.GZIMWY:^01\ZA#[36D=/.FH-X]1
G]c(9\gQ8SFEWW(;@2TMUT4KPX@@HOaLG=#_F7(SE0(18+ERbP:-SO)+d84.3U&Y
W7QA8@8aA)a4DNE.-T#;X-B9QNZ:_,:/W#Z95D^IZL@7FED8d=c7d6eIAf]^L;^Y
^N+-&@_,O8d+YQ6SR;WgSSO7eBa;:CID0-)X]QTG2I<CHeT+]6d_L4QIa>bD)W08
3[=QQ4(\>[@KN>fWD-.e#G8XgHe[9JSagXXCG\6D^#_&I\7X+ggLEe&gDG3SE3+<
J8,<g&M0W;(U#R;S7LFUX-@DRg7McZWRTU8+cLSDCJ.Q69@c,@/+SM[XXdL9@WMZ
Z@ZK>^LB/4U5T3UT<BY9f0+RO7+c9?2L<=BY_S6S4JfN42+8=4/(#++5)G_SbO3g
GGHMJKdO8(MW3YE:b/HLdE(@@/J@F@c-=<<3+-6KD>UMM:/O6&O?-VP#gDTDcV.O
^T)3>^df:OYDZTda#F0aG0\f2EKCOR#P5<[[eba[e&E),R+LB_d(\S,./H&8@ZE(
-b>L1@(J^QCdg7\IYK+;EVMBDV_#PgcUAO0e7M8#a+/7^B63JZY8CIT.S-E<+B?<
e6/WZdUAY6>-(CLB/e4CMf2:I3&[^=3-c^Cd(ND].7=5H71=-ECd7I[SP4__0H#=
S,MN\:6@OgYP;8X?cFcc6H-)]47ECYbQaU9OLG,6a22a[Cde#(\F^[DI72#V=Y>Z
OS5+db&JVLKC&06d7DI&&D;]D.^[&35fSc:TUe?QZ]P\5SOPdI>eCJ-ca;:fb?Hb
M(F@7Ub\[.YT7R[GFL=KX.X<^f5M_(7>>M>N^_1^_8Y#=2Sf6FY^EKgT^VQZP5_1
VdS>S5P\]#1a)UO,8H6OETg7TS0:eW?YB7T>&3Y-LZ^K95V#G3J<^BTOY,bD\;1f
f#F3:UZB=Q7BQ^(f/>VRYV9/E9ULg.-M2BHbPC3>7]/a-f:bfb8R)6e.Xbf.SU&3
S3,\bB96AMBY.T[>=;:69J#UcLTW9Y+30VTT[H3,R:-77SKPeJN9QL6-9+<=/_&Y
3Yd39T.+L>..2=4EC7Q7;HE7F3[-IY]59=:2fWGF]CSK=0##e[<9@>0.+6]WR/Z7
ce20Cg<X;#Ub/>TR6C+EK;L1H+QP<=;aXJU@VEQX.@<+M4=_)<Y7V,;/0Jg&[F;0
bPHe8--B9&=T;;gBG4T9SS<W/^M^(&<FLYV/@?YX;NC3F(;#GQ)EB6Ee#O2cfE85
CY-a8=M@Z41NKSTF]Jg#K4dE)I^?/8gTRPCaGC?BHD]AYD6KO#7c(Z8UW]SO_4L>
Ma.A,D?AICefJ:C\[gI@b2HP1T+efPc/0GWLPW8_,:a\4>g?VB.LZ\]QfOHB;7?#
Hg/H91\BF044(OOdg<Y^D&O@cC_PSP(M)c>L?&[GYce1VaOQ#dC]3]AY)NB+2^Cb
5[BTMW^D/ZMD/GE?=4DKY9D1\a1OC=S>Y@;,8B[^?1@6,8B/F\5]J3S]-H6T>N-B
(^?.4aZ^Ef2ZN[9/d3..A^d)deRH;O>.-b[c]g:8[229f,R&7&[,VI16RN0.G9&S
/&J:5f]((QVLV=aVQA]#Nfc=J#(Z2KIc&7d[g,9YVD/dI2XV.#L8<QK9cS^JHD=@
H1<_@G;P/e:9.6R\L)f0L+eg5VA2&VF+eOa(\DZ\KYU3G;SC9PR)A[NCH;>,)?/\
8gN\[L=BRS]eUQY3#@O2bMQ]GM:>LE#dJ\AgN@)]f&C6APA02\10:]TSdZ0P,C50
g:-8,UG8B(TBADGJ;BY4HHAYc\=303M9\a(/][](LE@2PF3?>c+J^ZKaeG)G61Y9
89CO5]:6#6dgE@66bE&VRLM]Re8[4^N9BP41E?0YLaUVJ1a6HO?fZ.D9gO^<W9fe
/aP#4U9Y\RLBLS/++O5ZM:d.1]SEM@A2F3BUaJAac&8@;,F)I\7IM(eO_b>KdC7_
:R&K7Fg/UR=WbCM4g+G1cD.=8.R+\NfF]gV(\D@cUR01DQ^dCJC+H[?bD\,7EYVf
DZ8J1d&;\_7(O:\=324-e2CB(Y9QA[=g0&(gbB8aU\GQG2O?)aZ7DC^.I0I4NdSB
)SUdK/g.Yc?U-M[<^#\F_JAL7f>3V&:U&1V;40=?<(a;)<,/G\GHOUP,5f6dEKJ3
#2=d6g#T]8bIAf.[RQYO<c\?NZ51b=A>7;9LOHD@b0)Adc<[4bB+]C8:aF,M&)^Y
Fa3-2d3QA2b?A,<8^/c0>[I@7^dO#72PBV:PQJWE20:UY+<I\851L8)<Bf+S_I_T
JYG(&O^[dJZS+-G?V5<2@gZY4R+R.\#;O;6bWaS4Q()OJ)K@Jb;E10EZ,9Z5^.1A
,6C_\a=JE9-a^3&9KKfI-Q8M0BJgFIY2;//aQ/KV9<[;4\DOS3HL1.fA#4aa.(FX
R__IM]-G-Q^g,7I16_792Wf)?HASL1XIL9(OS85&R(2DXB_W0d.S<8a-JeICZ&_;
@0_11W9g<[5CK?>#RgfCA0383)_G.I>gJcS41c18\@L0f5HS#.=9Ja@HP5(<eXFe
2H=0]dH2a+Y2.\UgJ-BC#1K6_W#].Kf-;;@8,,CbW9eV(C)(:\U5\D+](Ob(VDUV
#OI[8^H?bX?-URE@=V3AM#Y)K1P6U1R<C93OW>\VRIU,8JcC([),IgPTJ42T6)-O
R3=V]-;G3W=4Y=:C:7GJ6\3/P28EB=><;CMXQa&PL4?.DYGK:a;@IK:C1G(UdK8I
Z_JR,4\A@[7\?@dFT/FDa-Ue(9cETd]#gQ-Sc;=eTZC(6@\K:WAMc++5IEE^.OYA
52P-e<?JV-D?b;#)&=dN,LJ;CP[P9A4C[#a,74]2>0:;fTWf/7<bBeG5&f[S9B7L
&+@N[LMX4[:J=EIAA^dHfTATA4QgdHS9LHG82]@B?G&Z\5e1LJ6&I]B9Y8VJUUee
/E-?YP@feY]L93N4cSS,395c#fOG#X+Mca&-\&:I+Jc4gSM^I3IU9R^WQEL7RFGT
,#0;C.JKJ<_\A5=eNLFI[+_5U:1[9D4&QLJ([ZU]fG>,4UM18E1]5Y7c,g>)gJB/
O]ZW.^WRI)D@:NZQ<eKDT):;8?J=IV,JR7Y3)]X1e]<Z_;+0E)L@DQ26__+(^g&1
=IR5SM\US]33WVBBacWEa-Y,_8O-XN3:b=ZR0+-.DdgM-7I;O;:@M8ga;G3XX?<X
87MJDdV\d;M_0EN)@Ne\[_Yf_[M6HK[]QARdM_A)7OQH3(ZK.V[@OIBG8BB5M#b6
9B9eFJ/:,O_?M&3__Q(JBBW<RJXP>aW&;A2+;a\@8X\0>;RDUdYSL0>NYW-BS(1O
D8a(T+B^dQD>bZQ@M-V3E8&BN4LWNe\8AD7N?TT4N3#E(8>>+QISB=AHdW(7OeT&
H0<Fa[&^b&<VKEST9@1IXVO(WODS@2c8\P>V7IgF]TL#e[-S^bOA0X3S(3GZ#^J_
O#1PI=5PPMN14[RAJ)D:,&g.H.=f13f04g,gf9_7DMJS?/,OdF7N]/NF?=B:.\2&
fb1J=T,0OQMRaJ10LU9e3&ZTPXZH3PbeAgIQ#cA4(4^@SedPa2;>N+N^ce78+A(Y
:;J3;7TRBPR00&1GBCY27JGN8f527)e^9ZFF840T(<gcb_/_@Ke<HYfd,7H),.9[
Kd&:(eA.De_\b6:,(bGbT.FGg:If0a,O.[(R\?Bf_8K842?5D?_M/Te7H\8NBe0d
2.:/+=:9AHQZ8LcVG8dC/)66^3af&S<HBgE=_LP1<Ug/Sc5<P::J^C^^<(I2(TL5
Yd=]E()EGY=Ff^9S5=gKb>\Y60\SC>2c4U,HZ<P9]Ya&AQ675BVFgW-)>d\II2;:
F_P+b\@D7B;24M\7>>-<7U^-]IO.6M.0BeAO#?Z\VXW8EL,ea_^H(2=^4E9BFb-A
B(+B8YZ.:06&S[DDWM\[;P#LdCMZf&FW<&FH#X:_ScK<WI?F@SH&X/8\bX1Ga:RF
9ZgQUK,V1FRSdI-+7+I?\<MY?=7RQU^R]N)YSD3dU&&>M9g),g\2(CZUW]BHMFXb
b1ff<K@:FeG:,>8=1ZeC+c)0dHL9@E1:b/A;O8&I+K<PGQHD9d>g,<J3_P10+RUQ
bE>YBDTUHIS7EABB7Q/aU.OIcbT[DOFCS\@&,&S>fceK=^(1a_JOJ&1M>E4<b69)
G6aJ#Ca6Z1FC\[9(N?-2V=-7MGMUK-I#YLa7QSY#E1g91V?4P-fFS63H]F(6F1][
[fD1QLS2BfX^-/V?GI4g;<;LHMNLRI(8I)>&=Y;ScedLegVeSW([:=GX47>F8V\>
3YX;@<\KPQ@\M3dQIPNaa[&:G.)),@AMIKU:O/NSR:OYX\0U^,J80[AdUJ?@;N3L
9GPHBZ?]H_d^=?=W#??gHVg&VN[bV#L1LH8=0Nd79?&VVM#[](UY[>#AF?CH<g3A
]Rc5-=7[<b.^dIGSL&216d9Oc=F6I\cU#=+]X&:DM+X1ST8[EE,cXWbRBbK(#;5,
E\\4Ze(<DTU^8fB<TS#</:C^eRRG/MN31g.g2a&U3XReX3>eM_NP3/CYZY7-UW#,
K6FX(\#+E4WI?,f2bM-;U/C1+4@f06_T,0A^:GUZF@GaPI_Oa@g0M>;6NM2__S/B
b#U+D32^J1IVP0OCY8,0?+]3-;;T0BA>F(<=)RV[>?#P9AVdEW4,S?;87YEHgeZ@
&7L^=7E]eDL0eBd@4-;EeETE7f@JO<U.UZ3Y>EDY]N;gSgIU&Q#a(:Z:[W54/MAa
LBT7(S2a3fQ#c#IEG).28BM>BS77GCN9Bc]Q5ERT>>B7gb4fQ+dUI98_=M8gJHN;
B+59BVgCe,7@689gYfd,e;6XTD;U2;Y)e;8T9.XNA]7MSE3SS8.eAK:4[C1f5gL?
2_94c4X)=a?D@LGJKDd8:U7/OMFDHgE7L\B&M+682/MDe6P4-PS+JUXBJQBb_=E7
G^?RZN<Hb9&]/a&ZgQ[bD9W==2;@0eO?FZW9XYHd@;fCKFF2,Z->#QN1YVSKa:gX
d044XTYSKHW?H_<(H,fb[LceSF[MWUBF3IWQ(PJFA\;Z^SIFOSSTLYEfT:[KM_Ub
@<K3CP(d2R4U(cM]GXML_R2dQ^G+D;@[C6HNU@&LfbTECAI@PZL#7YTU[\1,ESRG
@Vd4FK>+#\/VUe]I.G+M9EJXTPMe#_P.eDHQ]AII+d-R.BW^XY=U[36GN@SPU&/(
O9fI+&IeZd(AM_KDYXLZXbDec)WZ34:O#,aT-TK4V6c;JRd:eFAP8+I:ba/]RTdY
LB_O#HHgC:)DW57@D2dZS19U-@Y1&AYH(3Z;]GSFgRc/6>K[#a\Y01F^V;I#^Vd3
dbg-M>S:;f/AM+Iee(EA,MC[0(9QK?)?DaO,c>A.)98<U45\U1IG_M;DPe?Q?aG?
Z.?^6O]CFM4,>9<JVISG:OE27cN),dT#.8-K=,Y1KfUfDQ+NDGC0G8IWELW_?\4G
cCL7gfaL(d]KT6(B5B2OO\fA)L#)LPOQSa&C.7D6(DIQ/K.cBPW&f&QTZfg^@:L1
>1dUEfE;+eF_F-8EPd5F@bN3D-;[f28DdMd7V^CSg@;R&T(<U9S2Mg4+?1aIZ/@Z
3C5_VA_YHLTfX[]-6QQ)T:gF2#7)Z.WDXA16FHO<Q)#VR3Ad6gcQ)#)56bFD<3+F
F-KD5cW<5M&d8?[e:T]XAfO:LBR\OAZ3_#S2T&95@+_-9=VRf#24.NRUY?L_(Y6b
d>^RVV-MgFR&OeMDPZR60)Y5P[VNIX.;2L\\D<M/3(d1QY?SKab.@81Y@UGaUR(5
=6AeL&e(0e1/6QN4HC=D89b)6aAB<dgfXE@0eJ\B&_^XgV(g)Q8[1K?I:-26O7Nf
]0(1<TgLIgSAWRG_C&3<cYRD[^O04FLYX]U62f./S3D4((4K?(5F:5;I5>14P/.]
LHX:?dD_KJY3.[7+.&QH8RWO#LMcL3UPLd3dEZd0cPL<6YO434SPY#?R9A18e.AL
.gZ-E#:N4Z4CcV=AS6QUWZW47;8R#,]WRP\_3d@J=&eEB\),5O1@bQfGF9FXNPKK
^Cb]78)SF0JI16O;\WYT-Sg-L@>fPb)D6>K04>6MgZ_?B>LBAK]D6Z_N58/W;:(<
BN(Z:Q,cEFTF9OW#U5PCZA^Y9/3@L<8_Fe8K)6YGA8\NJT/Z=A/(O0aT>IGO-f&0
\5Y6B8IGfdI0[)3gb9HU02fNPIGD6,SL^WJ,?eZY-3]-7-QIOA,R6B[Ze:E/ee:Y
.dJ_^L(J3JC^1FeB(_94F-SaDV#MU/D8GH3Kg89CSc1_cL])2eAX@+9<Z,g)TYG,
-8G=+J=9AL3AY)87N#)F,?LPbBb=KNgZZFIfeW=dV=/=HGF-&_+FFD_aX2McYUfV
(N4F:@<L:W5H5:9><VaIIWZT2#eQK1)&(V3/-J7fB>)1+ZVAe;KHd[OD5F]GZdO#
1_+Q=DA>5Uec:13<bF\Rc#,Q\KUE?MQ-URF(C4BAI.AMCT8>+5G985_3YV6[_C8Z
)8S9A]cEPdMXY5eRQQ9E<^5NBGcB9B9X>Cd(5B_9Z2S0/A4K&J^6EGTVL_c3F>bF
_Sb\2_+HP>7.MgXQ>ZIF0#[8T_>FQ)\^:008&V&ZdDBRZRZ2cGKPF)YX6./1BfgD
#/2,CR/QaYK33&fN[E=E)LA?H1C6H8b_(4\EX(A17S#=c-f)eEDQY/B2[d/fU;O.
c?^P6d#-bU9NTWOJ_)2&L&^#SFWTA#\U4Ca[91c.KRH)1d^FN0,.T/89WJW5S:Sg
WY]V]=T.QQ<3B)>6/PD/0>[;0Y^V>5&R?(?g53;?H/3XA^H>/c1c>?3;V3[2<(CD
@8T[-1XcALaRSCgd0G2Ee5e:.WA&&Y#fIcZ[FL[HH[aRA@MO\-->E9OF_[D#,d1#
49#+F6:PQ>&7E_#3?4.QQfJgNV@\\GZ3K,WgKN7f/LATb_B]\f8.1dMWTdReRc@O
d<]V=ETW/@]Rg-d^<64^^S,Vfa8\P89XPQ.9\,2V<T+X=Q?Pa7.WeXNaQARC,W2P
ZdOb<G8CGATf.>F<_6XXDN<ED?>c/4C4LF-;g;/g=#/81I=LGY2W]V<<GD1YWL&7
X@]RUW03P3aFNbVO:-[Ra5=G&3ID3,G.G/C:;dL->/O?A^PbgIVAQDfF5>aB>737
aL7ZCHJ>AQF47(=Z80VgVACO0+9g(6[@Fb1()YU1>)&P:#)F)):_Rb-IKL>VMO.f
:H2=c,4I@<2aLOHdLLPC]/C)1-IN2SELN9[>&+f2aRX;]MUBb?]^G1RX>2)g:=\1
dXb^OdM[J3_3RB4RUcWe1R,M_C2Pg[G/GY<5VAe-]a2/HJb=65gN\#SB</,E_fJB
SXgA^\HZ9-0\fc,ZF^B]AX0eR-+ES,P+.4c.Af]6GK3<RLMN_@?/]aDH)ZM6dR2]
M&?eZ3g/b<5SC,[_)Q,JB1#-X2QIP5gFFUMGX\H:HXDSXQV=0BgKL1X]KO<CJT4?
VUQ6WIc20.:PKcW378?(>O=<X(J89&BbdZB7Q(=[0F0f5N5)K11GCe9G-@M:I+A>
+A9G+,#2JTgHO.(RE)-PX2Q.\-]C=,F?1VNN+(XE53<PW02bf[_IdJI;JCQAc=FI
^OP=4M-T^Y^U\a6)](^GZB-NR]gE>a4F2CXXd3A(O35CG<S:PE<&ZbXd]bbP.T.<
@<#52FBU0D3ZO.W@e5//fC-Ze4ETcMSUd3=8@9C0C8+Z7O68TE@UU)9N/HP7YH07
;EX/>O2HW1]W#(N6FPB3C^KSRN)>HbLEIH]O@;KHK_6DKa^FAU]YQF\AB,VF;F2_
L=LD,e2W<EK1,O=YTeaeQ)D:H#R^0H#2A\-O<9=bR3Z=(].9W3#bB<4>[QR(Z96[
1<\//9YTQ7_/WA/I4BU@V2fY,+\A@EQKbHS;)8>AH29=C:^M;WKbHVRMCDCO3<=e
R)JGXW6?UO5/Vc(X3IQ=QVKC?BOeYVeW83<Ig^SV[K_0+[?2+ALd6XW28d:Y=V=@
3]c.\D4=_W9MO5]?5g+-3fV)de((#-HYCF1U^9fY1&bL3.>UcAJ[gG6GAH6fT,0A
K+0AFYgP,bKFg3HRaLbA__6^F8F_?;c+H8^a935VTT<=4SFg.+\G4HD8.AR1aI0.
7\R]7[D_7M@g#1IY9NEb@^1DR6O+TdIBP.IY&62RAY?BCMbQHd\b@\Pe]?MYHf1>
d+^.L\KA+=AYW0:BMURdCKE;WNUX\,@MRWN5T=,b:1KD6ca9AEE202FbHR9c0]<2
(G^LNbP\cJD9Ugf\6g=I1,HL&L3\HPYV73Q,XVJ<D?RN:+0VE0VGI_Bc[bTd83(@
e(/e2<-gdKGcgALB0VA:\?XNQ3HJ\-U@-ZRI^X8,_IL0bNLf0ISOFEc7;/,E:6[:
#[BQ5HM)&_=c:?JC;G?D5P&b4H(CB,N7A?E:dJ6I1&eI4=[4TCfTL]bZb44HQ7Gf
.4aTK2VB[>^.(X(W9^A]R6C,aRLb^/@T1;f0L8e=gZW^LRQYIT?7CRY[gLQIHDT[
Z;1[HZc6EcVK9<Pd)Q3YIM]_1S60a6UJ#-9CF=3Tc15R:1V&)_,\9\Z^WDfe7HMM
3<bG<ML:U.BOY]>3C3-(K\a)(TVa>6f(AM.7;)7/<AQRC3BK^gg;]<ZQB@,FZH.S
MP?dI)e>BCc_eG[-ASVG1F#-a:]#(U=29KQ0aXf<\K008B@((+UfCR&)gH_d;:(A
-@,QLJQSY_.a@B2]bA+D>9E#R\T^0>&345C2W\=K:@ASdMBW7<]H994R_SV4)CU:
2Ea^]<ef9(VK&d5]U[3NNd<c>a--a]]DC(TM]eG(1JFeB&/WLbSPSF8DW1&,f/UV
&AS+7QT#FaYH,Rg8f__2X0OI>c@\S0).7?TLJ&O1f-f-[0IW2WDJK\@D2C7QX.WH
a(8]UG4O)7@;G+Y&7_DKR=\CUDb[X&O==2[gd6R30,<6Pf.5SgUH?d:9_1R<N]<d
2Gc-0V<(T+C#5E,RQP:2IL.EZ#6YOG6ea45@:BX0\)J&AA0Hbb#:+V#]TWDR(/C<
>XSEfAa.Xa8:X96Zd5e^E;Q#Zge+g=/d^C[JQ#:P8VFN&Q-5>ABb/OGa].;,9B\Z
^9YMZS>,U98:9.OZDL.Z5LcIXDOFbJWO)JM4-9T:TR2CF.C4HI#<Q:,39.&.TNLM
O,CF@ebC:P-NE66A7B=2NM)+b;eR1(=]N[g)Z+D9MEB[8Z8OJZ2[(:OI3+>QD,aY
\N]_#]5KILD6?_#bAMVF7N83QBJf#><MV;B4+(HdH4]0T3:AV8VWW5QC]76P[LST
<UOA52(GA#L1ANJ-a/SCH\)B-/9W6=G(c#Z\:L0fXb]HXJ3E,:)DR<8a_DTOIQXd
4220#RDA_=DM.<K6\_4K,E@G@bb2L6Q^_VK;;7+E8b/BKgT\-V7<>fUG3a1BCaMY
Z?I[G?&+>V#<R6)C5d(6JdFCJJ<DbC39+LZ@L<6X(ICESMB.8(07@_WR(?EJU>-&
W#GALJdU?a^Ue^3@I7cY[D),9GE5g?[UPSQe&1,O,Y/7#]:?OJ1M_7-QE#aXE9+6
J6L]SW^@EU3=1YV=Kg2(Y(9S2<QH3^5W90,9LK7Z:J>9ZL^E+:BK/_2.#V#\HG(5
cF5+4f?aL]8.BHV#fIYT(>Q+.3(=bKQ,M@0#W)&L[a,U-??>0>GCgGAN@]M42GbJ
LJNCV)@bPZ.fF-I+55O<V:]c^?[.&/+DbETN.ZdZCHT#J.0cFc:(KK&G^&S[V1>;
eUG?5I6Jd1V7BU57K]dA\N,IZACM4##SeV=Q/Q_L4<C;GdB\dVdM=NKd+OO(J^)B
T<[(EAeV:BXf.?.b.Q_d@5Y9#\Y<cRJ(+RMQL\eX^#XXO66T_#gCdb&AS#1CWG0#
/<>0)M)Mga.^/2Q)bGHJ+[UO;&:YW]D>_#R4KQ7DB\Mb#\O#fgBENg7^S2S\GLF7
4#d0XcT;,L+8V8Y;#AS@I]&ZEJ4fJZW8>O<.>@W0aZ=WZ6I(Sd=gC=I=4BS.gSJ<
aF,SF<OWR44>(R=bW0CNN&BE<T0T,Wg=db(.GL;HK3IOX;<I[3_G<DV<6He.O(BH
[YVcM/ObU_UdPZ0.;?gXa2:7<,PNdR^FIY_WCBdMc/@-+ACT_64/COgI@\4S>9R]
L>^0+#I:>Ac2/3<7&G)#P?eP.+JI3;H05[9F0bV;_+T1EW27CSP=6NV,6=5;>3=d
Y^9b4f=_O@@]5NIYI?)E/CB<7<3F_K\A(@2+@5YLRE_Kc7c#4,:Y6LcJfW+<K+X-
T\5V?PeGF5L\\]?/cd[ULS1-G.8AFN4M+=X7BDe^^?Bc>>YaeeAOWe/+6G^VH44:
<>JM.Q(R8@a&)e6=LGJAagB]+(YWVVbTg>X),@\JC.XFR7GG@J)SZ,J:PU^c39#A
KHXT=[DINQg(,TE]4;BM4+fC_,G@#_gFXQ,PbgX,GK>QNX?-Dfa[Je?]4J><3Fd3
](HM3NAHKSQXd2P]@Vea.8;N<(#8>R(G)?97JG9(-DF=2WC98.4Af-,))P9Se.X&
\dH-\)KeL4+?7CF\W=-A5Q[=V[:__=AINJbEH>/O]Q.^ag>C#C#H4A-II?e?&_Dc
SIBdOHfIgC#^7MeB@OU(MEf7Lg^#VK,MdI[8B4^.]@:V:(<&</)T+RZ^R3:]^/:T
(5P6U\I5^1C/PV0XN4cb99P=52YA@\J,+72;eRK>BF;;^f#.dPb^=X#/QR;R(8UT
--Q<&:eF:<eDU4bLQJ1J]06cBY0O)Q,X.eW[>_a(2J>e0.FeX??:\^G@U/22:;,A
A(_R+@0@Sa=)?c6^<?UQ@P7S3cBL[a&a>>G_0VY8OU/62OJ(^K[g6ZV_6F+(Uc4-
c]02W1-6)beLe?a\2>E\U.>;W-ALeRDLf+R>cF,8H)+3CT#9M&Ta]73&CLL9/^ST
\2;O\V@Qe^]f^U3<,fFX2AQ\6fBfFLa18/?0XJI-;bY<^Q01\FXfY)S1;&0/&J27
K.<RZ_MDMH1YJ&Lc;S=)^8/A#L<cIQ4M0=c-&B_8_47T[@8&#F<g+-gLc6af+\eY
dGfE1.N:UU&W-CeZ;7K>.C\\/-QI^eT]CS&fXS+0)LQdd8JN7AN?<ZL0A?[aR:)Q
0@<O@8#U7cIO6,WDa^=EZ,L,#\?\5,=3FF^,4,GMfdgYR.IZdccYF/RK<^EYC?UW
#_Z-AEB4@\?VQS3&[A1eM@L@GDEA#A:Aa:cX(XNG,VaYfCfDI)KH-O=RP.G..8#Y
2f)JFE&HLN&O\=#5A.1Ug=QT^D]#SaJ&=R_[@16;6209fMKL.;O[F9QQ<c#N7F@Y
VbDH)<&^ISW?40YP[cLJ@NTW)C#3N<YA.VG6@1g_EYP(WW:1LH[8e6C\H5S>2]90
U#^]]R5^&(Se(d]f.FE7E3:6CcPTUC2Qgb]N0Nf>+2B>dFA&<#J5K_,4-c8/13\9
Vc)[.Q>1I3cO@-C3Y2G[A/;Yg.\5I6Hf<e#-dYGNMX)dRTY,Y\&BMc^,L^eU,Y8G
IJ5fA[\BR+:5O+A;#L<+OLHJ;RbVOfX(OgO_cUcBegbSdKY>0TV&&[BR&;,b/EN7
7GAD?YNPCB2LLb-O(9E&?J/(5?8WH;T+La[45abR#9c;_D7fZWMD,G:00f0ANTJH
;0>GeYY3TXCR--&UJCD^0d(L/G)4H[G32(SIU0=JP9C):_J0/f3]VYL]:[>g?;B3
;)#Ia<QG0?5,WQ;;,J@05(Tc0b<a9e(#4N(T8F1N9H7T:bJ0NG>ZP04^ZBF:g_[Z
#CR9JAE(-f4)]+DEG=Q[[CDfaG6K11VW?EC,Z25BBQ_Sg&O9AORa?;WVXSH4@_c+
Z;MbJ^MJ))05JE)D1O6;WbdX[>K]=?>?7)dL\IOUB@0T33J@V8US_1dT)=AZXX]b
4OX.NV<c&.ZIMP0IFHQLeIK>0[@Qbgc0Q0PE4c;MI6SK3-[85>fQKXB6A0/bN1@J
LOMd3Q3(]X5/FZ4A0ZXKbD0AH]7A<bgP\7g2aS+^J2e8cZ?9C_]G.[4SICC>F121
?VE[=X/&6/^)6gc@eN;#L<[D+T]UN\HReJ(Qgf.6Jb#OXbMKPT#dPA_\^5+^P>.Q
9-E&VH\g/J.Yc)Rb>(N0dZP&E3?)>L><?#.^4051>Bg3G4N;M&<(,GKg<OXGZ#\D
IGgdZ#LMFXXTKYL86@0=6A07Jd?g5/ZT-3I=I\TXR.+(f^F8efA.A=62[[:H]8QB
-F<dUPW@X8ed+IQ1<a/BXH(\S[Ua+<+#(Q]AC<IeDBP/FB7YH.GS.TA087(Y#EUM
UH,^;@8@bUdTZg3G>H>5NIfOJ2P][_MYCFX[WJL7J@1,5cC&3#F;J<c(#VV#H3ES
3LaF)>6;Q5#W;d/RS6WT]\H7^9QF=Q8gPe.:3JGKJ>dJH.a5Ra6(RI1VE#&?DNbA
P#V#54EUL+5R>](:\bXefM34BI^)(BMD7<_^-c#8D[]/:T(F]ZT7+Z(\Y&Ra[IIJ
V#+:TXeW#W1/?Ea-_D:VRX\g36Ab3MU(/W9g0A]Z.1F07=76(84KKOLFVaPVDZ15
11c8RJ4,OW[_(KJe<aN;gSI23ISGM4C9J/OXW/=GeM7X,Y8fFV^B692@^,58M6Ya
;>O];8W_NQ5^:S-E>^EN,TXKd:CVaY5fIN0/;O5FW8O,B1#D3BLd_X]Ud]]c,]UX
LVW@::/=QIGKUQ[dFVBBRSF&&T21_C;X#SA8Q0U)U3LZK)JT).Q;_>(,ZBFQa4J@
KfD\B<W:dD=C32/?dQP1HAV@AJLR(2HfZ51afPTO@D;@+P0T,^+7]0HG^:fSKC\K
>=.)MgcF_Ybc^:I\V-;<F1GVG7NMKX4(GOKRdYWg,Ec+3?-6[KPgg?8XGGd/b>gZ
7W-G;&(b5:/?L:PK6HG>0<c<eZICaJYY/RfMR,ME,03CNWg?&eX;\\@IJb>S2[AG
6LOf4df@UST>WGWTf/FPURJ&<#1<)C2+Va:T5eO2RB\21X6(1J6-=N,)WIIf@GJf
Q;b#R+XR7OMM13^02J2KDA6:0XcAV_F]\,eZ8QC00?4Af3<8H5<Z^F],=QBUGC/M
V_cROCRaM980M@GaU^,\CXe9V10BQ;5-dRbZ6KEX)HKGHgUY>[Qc-@BSF6U-BL+G
cIH:-:f/K-62SWKFEf]TBA6\bd_I&WbWb6UPD>A9ONO,N-X^Y.F#QfFG#gC\18T1
2#5c\bH^V)^c_Z1,6253NQe]GZe<\Z/#OFX(3H4#CL;>QRX0J]APR6/X)6X;YfBH
I47d[R;?Rd-Gc(7?OC.I//f^EM?d=PC4aV)_Z?Rf#M)3@KXWc-B7E)>49]c+(QV4
S1490TF4L3g,W]DaI<^)3[6HSg>gWBT@6d_:=7#<d.c7]G+d6A)X&E<9<>gF35fG
d^g#G/)D+-7K<4.B4Pf8N[CH7a:0dLC,gZ-+RSX82GT5-@H,7[9X_^IKE(S.SN7&
4bB2c</:M-<bT>@E,fd^7C]=/F\)d-(Mca;EdW2]>&IP,I.f[T;IE827>97TMe?Q
7AENAO2.9]=dQ)E;ZaS+:f6=VFBG:RPd^T-eS3X<]dFM7)R,@/6+,BNZe[J0VQTX
\dU[]IQP=T15W0@5;,3L&E/1^0-R]4f]5Tb(.IU[XQGefRcO?F+O=#b2:17:ILQ^
S&^SeL@4G.<S#b)[9>2U6/G=c3H2B/bI\E[g3f+U/4fbdTDbeVSb[I:&Y:IL^30e
][LXZ<:Z6U;3QH6(N?=E)(KJ#^OcZ[dKMTb1,.RA]+eXYfZO7/9d]JBEWZ\<57D4
79QDP@I3b8@Ba,0F2OWN[dT1aIFPUM5fEJ7a\P3#+dg_H30JT\KL6Gd:W[CgQ+YD
9=Y&]b9AfH/ZPTHHU=M\4TKg4]RSOB5bS8K_X]DN<LPg&_52:YDF1G.QU7b_\f=:
C]EVNdV=RCdV6,.,_&44Hb?[a8E),J3W<>LTW>8TMYV/b,]aWd::6^Yg,fWTBLc;
((VN>g0:ANfOUM=+d8?PJf2@JRb>#\?/bBTbbB1.E#RL^\BD1U#W2G7f255.J^c\
OW-5;8g=ZB9Z3UL1AS^50\)O-g;-LY(0]<EfS7_Mf<T);&0:QPcHgXAD/dA7:+=d
c/14>85]KJ^+?b=-9&(3S6K0?SDW/+f/\E.9-KFS=3/^ZdOG,d0,YEg?14YHdb(4
R1/D?D5+eWFf.7&/G(V](.S,2DVSYW4bb_Ne.\@H^SOW@O0bd7JW^fgAG\Fd(^HD
3MUNSCRNMU1beCFd5I9-?b-1JfNK73=C,^2Vc?daLTSS6.E:@E)N#UCXbB?\Q6X8
3/02S#7a9RG&]gb0)^0C;P(4BVa4L_a5U-&R6A?&:W4B#E^-LUd@)R+ZP+ZbESag
^22HG5aFH@SC;HSeM8f9a?N72f.V14>\R82S_#)F6KD9X7?bc@3??Ca6EKO=3.=9
YW#E6;.>eAYK[/DBT5LO9Q+YZVd2cZ_;:N_#f#.ZV<R,427XB(BVF[f@@SaR6/)V
,[5Q?3dFG;9fc.T7IO@IG],3(_VMC58KA^2Y4G_&^._DZ?U74b2A^AbF]RfS(9:(
B?Y1bdA/Y2]TNJ7Z(71=ER2OUdC0E]>G/L_;89Ug-e>>9;+:IOCPM+)>?>V:bM.^
b].Z2\7?[1,G:U=TM7(&PgaP0aC(I5\^5/KX0/1D[@;.g@RQ/-/\^HaW(HXTKg3W
XS]77[6]^g4((eb]1_6@Y?XQbF6>X)HJg+S/FGS=\8b^&V-N_#EDM=1BS[@;1dbX
(8G5bOEB)+H-gL<LS<=aLV[(eI9/,Mb7UAG]Tgc#:<ATC)S@Qa1#Q_W+ETJN,fMG
g8A\JOAJb+XF(#aDa^X2O?H@G>74+1Xd4W?We,)O8ae\c54O@c9LV1;&5a.@#QLX
0\ecW;0@=&.VU@fYH^[6VKZXWdDBY6RSfA_[9:/#7\/HZ9H7cL=4C#>7FF[.M?6.
(2+29c]NA@X1R:\1Y=J4PJKOD[I2_B[K/J\3Dc<ZH&@CM],I8:A:LT2=fN:RO;Hc
Q:OTfD3aL]>T8fLM<Wg]JH#&Z4)O2GLN2UT+CJ#b7(XF@?XXVP5D4L_?.CS2Q,DW
D(]5+a:NM]URMXI081.T[L<a^F[0&=-6&QX5E&(_SYb/cXW4H&)=eCNI#JY9,#->
-((8@W&d[K\.UTe(L+EX<gcP=Y_?Ig861-&8\/C#3]d0.cfTU>58SZae4=82O<2B
38gcR9HC\R:_VF.&6IJVWNgS_6.-cK)RF:B0LgbdQ-P)ZE#O@642[LaQ^UEB]8PX
#4]P59g-9T=4ZFYfg-RJdcDU7N=8G#:=Q8R)Od#TU&9Y2fEZ^C^a^3<>C-e0+HYU
;Je663,@Qf&:9JQJ[.S<O<54+K#eZC37>R/f/e?bOGQcg:NSOR05TJWJd6/_H#3d
fEMS+2GfQS.Sbb1_&PDELQ#KLFcM<FEc2PTK&Hb;81SRDVR=KE>+8QU[4KNDVegL
QCeAL:5,Oc0-SY9L4D3bY_W]1IcN9_1aRc5\JDbW2f:KHL)1AfgT17ISXScLWECQ
3gU)IQ@:RDL5<Q1Ob4_c1,[Db.UTdD?Q05bV&+f:V=BT/G^=ZY)5+(#8)?EacaV+
EO/]E\NWbKEH<ACG1OUZ0@,Md3XLSG8N)..HDCK).=4/RLg[H]2?]G05eI9YXGGI
dL1_21@^7CA+UJZV9f\-PO)[7.,9YWc05b9=beCASI34bJfGDYA0S=6=&35Rb?9/
)\4G[C,eL[MC:_d^,43..bQ1,Y8?GS:6P+c_[O>W[&eH-EE)RVU_A^#eL8fR@aYH
=L38<.T5d;9YZN7@GSX09<L49\/Ma)J.6:Ba/6I>=8<\Y+@)),aS7Lg]fLV4D<ZM
S(FSGZ0I^:CKEZ?-IV4C(M2c0=G&H<=)&.LW26K=C(Lg;2AR:B+aFC&/g;KX5KI3
5?=ga8M-9UZH1@LT46U;.P5FTN-XEEA:#UWEZ\2NF\?:-]-=9HV?ZLGO>?<20CUC
+&DRN#RF-T9FB6+_e5Y->MALAUC[H&EE1cS;0L2VYOa4?)Jf4aGH9.C43\E4+M&]
(-,M(X9gX<=NIPQf;)J]ZXBKME<CGSfBa9DF>\PQLK06^=9?RL)DL5FUZT(K:/>E
2]a^:][-Q93WbK/Y(4&&=V3IbDD7#)+gN(dTMM<b0Z]2L>)VcNTE-Jfa+2[O2J4L
>LBZa:^FDbf(5ISLDF)RP7-g._QL(;a?7.H3P>/T9C3,A14G<H\X>?55JTT7Z^c+
J>11P1:XR,-#-3D4e8C<:^;T;G3<A(5.6---N0OT\Vg(PXK/fZeJ]:Q\f==S,FO1
)]NDCW6Ced&53WUIB_1(bCfG;?@Of.Cdb1[S?A&)O&W14?R91V74GI@KFD0LTDN5
061_U+-bB788FAaf0g;IYYbF_\6XFGgcHLK:WYb,V5d#S4POc=0SL9&K1V&9QO9[
g(\(UcLXcY)4P7#aQP:)-Z]7dbXX]7W75cSRW5[FND_c=N7.?SC3MRVU=gIgC&Fe
fPC,Df+<&8aGB_I]FMYCHS&45SW&D:1&bS6)^WBa+EL9_.CQIFP6UFUDCF6P#V=F
[;X>_1b8U1W[FGDMB6.^[Z/LGW3E,18aSIBe&G82aVDGR.g4U(09a5-6Y):R)U8E
Y(0Z&,S]eVX[)C,(DNLG734+#QgV&@L)M,>:]8^J4,eWQe9L[IF6?4D0Ee?#gOJa
?2R4:V15[-6#AcQG)EW#OFQR8CVfA62=^2JWb):cXIDA-e+LJFaA9)^MZ,9EB=RV
gDJ5Z2^eRI8e]O.Z[-gJ84,adbYDL\[/TJfW8O[P4KWe_Z#70c[EBG+X1#TLV-:P
LBSC:eE7(.2SMGC4I9SgOAG,3<\,a]0d8<XTeAPF0A\3-@Z>]L3Nc#a:P>,g_bOX
M4MR>fU<;Id5:TYQX\#VPHgUGUBb5Z_?fH7E-Z@O@F0U3cQH+2\D54g7CYdfJd>b
X(a:#b/X@f+)E5X)JVF<<c)2JLS)2.8^4&/J-BW0BKJ))<)0f.f0R_4d^<X19F9Y
6Q/.AObSIaD\=NHLL6GdN+H4=B\(+D^PA1-[C::G/G6[_KcNgM3AQJ_K.>:]E]@\
^Z/_U:G?RCH1GXV86U1?FI]UL&6gDg\gd<FG,eJF->&=B1eVR:-dG[LIeFeVU?/V
R>^>@1Cg3:gbYb(U8(X+EGA6>9BfV(-K8Y_NJ3?WP+=Hb?D.4YMN5CG1D7&I=^a\
)7V3<75S>a1.J4]&09_U_3c,0#&W2)B42_Z]U,U7L(O7#+15c#Xb;D(BUZK5,)6;
(I@OS6]7J]4D#0XRXU2_;bfbUAQ>@Qb1:/#O#-I^f8?#?0;bVUR^36Q7-+80U[g>
,NEC2ILY:HV3=759F,AXZB(YPV6I]4J/YYgZc7bd;B^,5M?=BJDc7@C1&9BK_Q)[
43?O<=/-0e5WHLF9EV>1/-AB73CgG]TD5A;-H).3:+##b.9BV;XV2U+WR8@5QYPW
a9[;GEE/[AbR/2H=\Q[;5U[]4:&97:DA^^#LI(?54260-LbReZT4aO^N0g<FA,LK
IBT7F>X@5CY,(Y@<3B_=L1cJ@QFYWPV97294Af;fc@V(b,&PM@/(f^[a+>^;M@SX
ZcTZ&R+VK;TKLEX1cL_),LXGD^>WS=U33E&SNF1((Q<;>[dL12<[I1Af5:0<dFJ=
[8cSgQRN&,+GN<\7+fdZL(-b)-BgD:b_81?PZ0LE?S6\/,=aP<<#Z:B0,5_Eba^]
96;,+5ZLG\.8/BHA=\;]L+AJLVC0C6KQXaMO5W]UbZ42:-RWReV?;f0aLcK3DB)M
;]d;=1#OTA0W?SJ_fc^(PBI=TF&=fL;Z\b:AaV?&55NJL+@8HMTKFc,TaL4I8A4D
b.AP1&dZBLA<KMFVXe&]EGUe91=-6,T568YdMd3-c3^,GKN;UZ42JA8?JS0-MbCO
T2/SXY27b#U9H<ZS/50MO9aZN].N]^9T,?SIg?c.CZa42S[2RG-.[EA,<AX,CYg=
WB^<;Z[^8NL+dNM:Q<_5(+dA47]Y2#]N@\Z\_X^QdMVFe5Y4?JcI5T<BPWO#8RSS
3Y@K^Kg(fK];.:dfC@=CGYQSM)Y+?M0[?48K,VPS>(I--T:T1_4-.\Ta,M,7R,Hb
\0)dZEcR@&3EX.02.?WN_FIKG?+8PV>=5V>4.fe#J8&],DGQ:QV4QYgS_\IRD@CJ
\25<2/_CDb,a/QMB@DML.D3M?_658K\&Uc@12)1X]9O/Qd3ZT+F)#.ZI=/DK:c;0
Cb;c95<BA=WfS3Uc027N&][EFRHF-1X9L(\+)(@[>N^9@23e<08@gWUNeTS(/G.Y
W:(b@:ge,UH^a:6V,X++P0BSRXAM^3Ee,M-M#)D^;>XT2L\,N7:S7#_<FW0ZP=0a
cdD/?Sb<3&?K-YQT@f)]dBEUeYRPO+6#bA2>B7U<29>M7<X4JbN,,/59e0[V8O<d
J(FWf3DIA9KK0.?7S&eTHbLKa,,agX2,UebCRZC^^)KTDBA-7B-a4?MZ&(Y6:UF=
E,B,gY6=WTI8H_9XAF.fZ1G9VBY0237&(VZ:?G1-AL+]<V@N]_EY0N,eARV0JW9;
XE@:)NGF4:O?_;@gDD1O21Y\Q1D_O+Yc<gVLb=:QdX[.KJ3YHX98KKgK2VCZFQOe
QJ=e:5JZRRRD;eOY-XNQb/JC<O0D4_>Y:\c3LT,TNX5=\_19VB6UM0gX)#KB]LdA
G48ESS/5S00\V?5,/841HR<T0=.1@(KJ^:^#AOeTF)J^__b)+b#&UAaQgQKKcef/
\0C?EWW=^]_4.NV?2T.EB@dNL#7=0V2QB;=L4P7/:>dFHQ(PA=^^8J6(U7;Nf69K
8^#S6F(/:6ZDJ18,,P-c/P&X5ZHK]3^/OL\^^,PKKMJFISLe2GMZ;#1@F^c^#K;G
V?<JJ<9Q\RZf/UfW:)5e^9TAENJ^79aS/fba:]JZXD@W9[5OJW[[M1BD5:(+2N0Z
3@Sf)NV6.6/7=>F0F>SNS&&:^=cB,?A7QQUGMOZ6c8T-JgNSDJ)B,;VM.)SRGWQZ
D015QT9MX=[4TG+C0ZDL)X.^Y:Xf\I6VTEQ+MTY8:2^JB.-DR[85FC)(UHWKKEd)
X1(Y\g@7:8cU+JaCJ#>cARBHKT2F)U1g.HK-Df8X:>Lfc<5G#?HdA>QRGJAed:_\
_W9ceg>Cg[g=OZ\gO@/N,FF[+C@.3c[/KI,;BZ,CA>:?VFWF,eRR-8@&YA#NO__c
0GIb(Q9FcZ+0)-9GfY:,F:3@.\JgO_9S/QfBUV\WgaMG6]c0F]N\Q;)Ed,N6J&F#
N9L9[U=>gWd.@g5.@8&g2a(^/<9gD8,)(C.X_d>=S]VW#D25:6-FfA=aKX)Q?d0U
8KcN(3L5UfD4T1G^8.\NE@[=;W1MEUfVP:DgS9XJ;cH0.VMAKOK..SX_=UgJ_:8H
1N]d]Rc\8;-<S+b&?,?Fg]M^(Ma6bgZ,J=,N<-BJWAe_9A4g0-MaFe\CCBMa,Z3W
dK)W238UT\W71fC#c\>DHPdM6GGR5WJc.4fN.>).5M8GPVX>f&fRbYBeQ3/-(1Aa
WT1CRMD4-Yde88^g9L)RbNa]-N^R9&K4Bbd?:/c+^YQ4\V6K:d[>,WMXPbLP\P?]
<?P.Y.K02/?898ZJ._8g;^@:][R3#8X9EBW/:3QB8gF7+P@HNL;G-eHURP]<9IBD
@F^e:YB-Ce2dD:RY3V+(R377160RW-[B1KdEGNG1AETDXW\O_B9=M>_(E[JDGRB6
cMX;3&dWKT=.d]T2K6S@&TTPR35f1Hg.4///-J0]2_KYHg9XX:=Dg3+F=Q&?X[c;
?bM[af;L#=feFK-]Y&2b01T1&f7>_YMD\RAJ5&6<Pe497&<NF6?f)NB]^bbXEKQF
I@0SYfSR<J_,Q[99&1gcITE8)NccHf+;2SSNFWc26Ac)B?-?Sd_aMcaadI-#Ha]Q
V2GE4PM=8B25^a1B<3Y-SC&TC;\:SLA:]G?3OLDe4/<45cXT-fN8SS#4FEB?[XS3
Ya;g7U8^[(Q7RL(b,Ff-1=;35b6L[-7YNOLa,Y-:g=;PAT#9<<8bAU>CH/(YQ:9@
TI3?DQe@g2CfbdNfd4<<]X((78GL,]_dg>F;@Wg7DSNU:VI<K?Z;F>T=,N[>>f->
X08?549][FT.(6/JTKUW\05]ZCNe<N6,;f5@S5>e5DQ(gF>+7Ac/I-87^I4>If4J
FF)H7YFD><4L,W1Z>-EdEOV5RCFWG_P&Q/cS1RHLE3O9D34=S(,-4Q(^Z\2ZM2-?
CS?1L(,U7][-I.dg4DEWf<e&VKQJ?f@<aCLV:,J2d@_Z?S@W6)^=a4_?T;<+WI.N
X=)NQ+gR_TE(.?a<A&3OYW\,.=a^)_f&LWdfFgJEV-I.H8B-3<Zf#K3<X1?<DABP
K4WDM+CK?4@-dMEH[J6)d[N3U3]+gNJREWZ#U8(_CbP0=[/DfEdb9G8G6]E3X3.L
\HM(Z,/A3dC-O3eKOF&K.KA9cD_18:(^:).8,LGNMd4TX(+d:O+/#=+VJ0b43UJ[
Bf&eX99G.AHUHX>E=JX]]HOAPQ&R.&Tec3F80;;GCgSTU=Ig_+XB5G(#Fa35(bFR
>eQ7&XgQeb;<M0Z2RdcA7^1_aEZ,J=#Z^:X3EN4f[D+ce)+d.@3(NK7\1@C84Vg)
2dXD1bZ<g/OXS<IGH.TYb^aY;[)^C-JQbGX6eN=5;QeA,dWE4K,-CO=CTVT+eX^a
(/61(0>&70FbWRQgX0[C98KI;+?/#Q;G0SYPY9aB^e(_<e8[8THXBGbRd5E]:FXG
:W9V+AI4Y:,f/W[Z;.gA0dI4[>Cg1/aRE0+;)QT-BL)>ZC4b^[[?E?CMd\TXGKE^
WT+:B9Z&e;&-79JM0DN^)/Ha9>USZgC@#6:@&YG6W4+I89+QN>K)F0:=;?(4T0Wg
K8@GIWcZ[:G5W+XB[3Q_M7-]a?e<f5Q_-CaC;.SVUPeV0TAID7:_d_&-We6#/A&9
Y2E]#7d8e9&)QHK,OFNKXTgVKLIS+dLAfXd/IdR4;ZRQ4X_E5FMg\;.;KP-CA2KY
?H-L826N[JXBM(P?R+D4HBX])I#dIObQV-C\9G\Va4f.7_g,-GEE)a]#=LO9f#/;
6gF>TcPd<(AB2GX4F@1[Dd=;.?Q^?;(e1Y#).H^D;J76S)\@UR_/U;SVSZ@&^.U1
2b]XFHIQR7bKe27G<DY7ISaaM7#/WSZE-dZ8b[:ERKfE6)Z\Nf[U2fK?18HMWFAK
<6cG9W^<g5FG3>KGY7)UKY1.1WW2\WD:daf+0Y#;8ceE6Z1>e=\O.XL\C0fY:4X;
b.32:\1DUe5C990M\:Q=S9RLa<c\eTZU9G=H.bASKD0Yb-B2EK;]&-0(\E:QD#N4
;-(f,1JXCY?<fW+EML[_4W/&fFD/dU,#;#_HP8X7ZW-_B2^(=IM/##U]Zf?BTeGC
/?\GDY6TbWF7R6gTTQR>9GLGXLM7@EK0/L5+6R>Rfe=2^JUMTP,HCECKZbK4<?XW
QTJ<e0,W8^KPLGTXDRG=P^CNK4_7ZQ_K.<?:EG9VW5&NcLM(aCPOgOF&C+E?>;E:
d:1fa#IXR&.U>@84cMOT9L^4ZNEZN5.G9>.V;K.aB?EYD[(1)F44_2_6dBIPDJX+
L<)eRAbWK-#8Y]D4_)9<K6XC?G]KZ&7B2G\GL&cDB6=4R3[)cZ<UI_./9GFM9,CZ
^3RQf?Ec(e@YdD]ZS)/?#UY-1.SFW7(Ac6MTIOI&N&;+6,:YH&F]5GJFd]5Q=J3M
VP7[DCSWGK[LPI9>TTNN=Bg9E0GJ2&M:1a\-OVG\bRY#15gf=]@K=DL^@a^#@7a;
b6THWW:>QTUS_8^-(?3DXJA<11>#\XOcRb3.-DaJ&c8@IbNE4^E0K//Y@G&\KS3@
N:WG/LN-&^EEFU2M4E8c&)4CdN^DC5fXfWBUNQE]\][=X^f&4>C4R=3]f(@W5d1D
#<O,9cVM9Z::Q?.^(/3S@.NW]IXSa3#PV(8>ZHgKdH67&V[bBLK(@(2_W[-G0>WG
/1IcUIU?=[MU(ceBga15g^23^L;5;4E&^VDS[L)9HfbV;KWY3.&H^G8MaMda2O/U
8DZ[-Ee2eA)@^JA1d2F)NcID[XR;^+5b<>>VNfKeQSR[Z?-F(_(f0E97A)5B0\UX
5I1,VHT?GDE7d4<Z,8e1F#H<MO]-DKVF3bF,DL>+fU;8Z^-SB>c?E(ddN.5P/Na\
>af81,8&U3[KV@gSa^NN3gNfE;bNL(][_KaeXb(WSdAcLSf1#FcaY)X?/@dZ[4&+
469(6/?PKXJ+Xe,..:5GO)G.Y1]#7SK)cN38@8GCLATg];JCc/ZCX;C937b<)F[R
/0ePQL2ea1,N_fWaPP+-_/)7]WYa-(H;R(]f+Wc;0]A?Bg]IXaE(/[MZL3[RUP4U
6F?Z;B]=[-YgEOd\Y?PMH@@RFPT0-;#RCC3Z2XN_gMQV]LfOb1PN9H8@C/\\c+H[
.[[ZKF(HFUAb=4R[PQ#gRg;CN54E\=-196\C\C@_IAJP_QBa+J9JB;5.(FO/[D]>
\Xb>aH>CC^g;La(F8_McZP/;[:D6FDCNB<a#cZF>N)S5#B^gM85<0S(@bA8HDL?M
>/2XREJde]0WAZ^\JEW<G[#T4Bba2?/[&?[.G2FK<WEKXg/0GQLC0^C4M57;&4E]
fgMP&&NH7MHQMMee+1CULLJ&HMKUB<8KTUH<OJB_\[ZB=@&gca:V,3<=#=I-R7A0
KR5VP-33LV1bS?A:C^V#YP@b=KcT0W)f<:0ROY)()M]>K4I4WKFB0\6?aSVG=JJF
S[H:\-)M52C04f;Wge-KT4_SOdgB>H&NHf&DQP4;MXUUEHbHEe4O8R>acc1b/E(M
g9;QI;M:.;eQ60^@4YY5_^c/0NV?a@eV6@BHF7fUMaDI,@4(WbCKK0Z.^J&c=V(;
V[:WdIaAZO2c+A_gG6XD3T_6Y+9/=N40IN\=5W.V=fK9NJ?/;;S9H3#D/V)UI(d4
FD6FY\;YLPABa9eBT_<d_;1-M]e\E9.F7g&&gfA&VHR=@^0<A<A;a<g(OG=M]S>[
TYe##0TZNW=L#UA&G/CL+=9)Y<e:+6+,TLZ-PN:a5(#^1d/CKf>TZO:?2,;JT<3K
C85,9MfCX23WeB/\8)T2^gU^\UK:4bJg@T?beM8^W],GD[d+bNgTVbFabL7c>UZB
6-6&KY<dZO<3X=?U<M@Q8f7\;AL,YeE;O+;;g6G][ZeWe0NN#IJ5P1/Pgd(X;W\L
M_EgCW+_IX_QOPJBK0gPGAW?/MeH&:F7O@_K9);fXME@ZUMPRGQQ3B:20B2.Ig>T
3M>E^XXZ]JGBU5W#_/^GgL]L@#\2LID0LJ=@_R5gBP)EVeOV4N-B\Pc[?ZBK&KQX
-b6e<?2\U)aH.fPS][#PW8WYBE7P.:PD;PD8S3)@#V#JH<V5R[R.;RR^R=cIB#Cb
X=Z@7X;@dA1bM(&c-<[T&]\;P4A5ZegMIIE+/\YgC]F<LGWRVV7,097)E(:W7+a>
9[6+cb[DeF4L#)1N72]:;S@E,<aU;FS@?UdFG4H2:UA:=?J=S#bSe)IXA#I0:Ud5
\@J.I.2WZ>#^K4db>)ZS1C[JKV3_dC>56Ug0fQH#3TT+OF@4e,Y09CVJTIV_&6^=
C_T:<P>6cS;]VN5g3MJ\)e]^1:3Ug#LgLaRg#REaM7W4A:@[DAJ@6aRgD53I;?R]
C@YN\(4[>fc&#HP5fRDd+4BW=VfYI>HYZDfQ+L7aL8AAfP)g+-DEHQ/[JQRe-YIY
^F5d,bT\ZO4/fc9WH4Y#,QL[5(>\=^NN@(9Scc5aLTII#HDVK@FG_=B8_9cZ/KN4
.DR,PL1aG7>-=03)a[9B:]A>>_@BQ)>HL^+A>&)=Ge\,T.&?>EMa4MB[VWD\YT2R
;8Q(@3\MPTR>>-[5e\b&].HJ3_LK\<R>S.#^AS&b2\R?-1>LC]c#0;/d:VJ6KD(c
5g)&fS<N5U-f[^K(>R4?eNY;(5Z-:6eP?M&/_//,\;dEBg&d.eE&+0>C.Ig0I_9-
BOWLH8=J&8OZVg(\4MC0#7T8BR?ZL<31g+/CSJ7[&/P,I?Y_B]K;ZT6M62b9e0KX
:0J47Ng.M+M-DP.328V(V(RLVUVdb?ege>56EZIMR/5)bdFPg+1/[&Fa4(Hf.4<b
T)5b)>LEKV?XU+bDH=9Y6T8/;#2N)E5MP=;KWbK&X+F3gc1?/]N\FY:d8<=#582]
=H#FA+<4[7_a14=@9E_8=7b2g3#]+-^(S3W4/(2KC5X_a<1B?9P(Kdb8[e&VH-[2
_U5D.V_Z/[QJPGba1g-@HNA,K@J5NI<\N[aB0FZ#8VT+#WK[KP;#)Jd33&WB9_M6
593X5B97RJ]7^<A1J<J/5XaHGWU@J7/9B>:UJ,7S=b1T3H5Y;M-QR+=/ORBBNgP5
gC&VEI=KdL9Y,bGU5ZUU.b<eWeVYVc=Rd56cM&8^fYT8)+3MZ0[J8/?_HL+06K0?
_\\21U^M9O<cCgX#Q)Ba,K9Cd;V8>H0SC>[KEP/4faFfOIU,BWe_^+1.M5gMKd3=
)XTYa6@52R2Z?fVe@Y[VbC;J:QTLK7[PM4b(dYD(_dIb,CFD9N_ZA(9UPe7ZCL^+
?-@:X1WVDbPK@TAOKU0W/SYEBG;/f>aV@)K/Aaf?&RG\-C5M&eL;--9AAG10F[^_
@H8=f>:29EM)&e0LSLeZ;#\O,gd:^<KS@R<A&1U<;)d:JIe1SS>0=(<RUb+a8V/>
>XdX?3IZg]T)\8\CYY6K\T19J)98D&JG6f43UXaX&+;J)]g-;E)1F6.5T>aY^8<)
X^X>L+bR95I/,4^ca2/<0^C:W[3FbKU,B5(fEZ9\UdR&3?4H?SM655#J==O,fK5D
g/+.^7g4C;FRVPgRW;]E@#P#M1G:UYJ^0/1]SC3FG,c1^./RgKH9A+4a8c[HQ4c_
<.)GOVH7Z6V=S(WS8Cg-S\L-+TY)+OWVWT/>c]UKbTdS&G-^FO2N)7:^&:e6<R,/
aNW.<7#g.3W&e\7=EHKA;&X#DJgGH_D[YBRM9.75I_4]]/UTbSdH9JS@QY5@),g0
He2ILMcZ_^@HZ^L#Ra8GV,?ee87-=U7A?H>^\V?FVP#41gX<:T>XJcd]G&TYL.<1
]1eff9MZ6[WI#E&?30@V#UIGJ,8fHN0a8MW_6<ggWI);D?U>T,G8K+65>>0SOfVO
a-aY7STZ/LA\4>LNJYFb:#W,TO>OG,&U3SFW:Z/F/4Le9YJR8424[^f3UT=KBbDH
.C\R#Z>;BW:]HF+NLE)f_<@EV#H50I[7Q:\[H&HG8CIgf_D@+W);Se?g0P=&RD1I
E?U4@[7P39YF0@f?eSAgK3efdM2(aGCa)/161ZO13O\2>7^)ODZ]=\]ZMfY8QKPa
HBS&(8O1)e_S;5.P@&:9X8MMe1GHUJ0C+#^YE6Z,UX^C5eXNeV0fZJ<^b[QF4]H)
N7dCV+K7Y>@ILLK.UC&=WZdC(..\IU&Q^I#B4Pg#@(Ka@)_Bg19gcU,?EOMYHJI3
?^PEZEDObH3GH:[E-6SDTAc;fWX+Yc&(/K^.>F4d9>K8Y@BD2GPXT8I60LU-5gWJ
7?SRTaR??cTZ?eHCSF4aW>Nf\AX9eLAWbQN7SJ3DHJO>YfcZ5V@]:b?09OQ:CX;:
XZK?c@^bP\CG>B:[.F;b)XTV-fV_IbA,<JA=b>?DYR(U20B6=68KN0P2=29]a2RU
+8d5<Q^9]@A1-F^UH])I<X6\;IfL6,KW/5@\BLD&XVe>RU//)E>TfBCOO7f\HP_-
&g/(@B1+C4,51K(,A:3YV5Z_@Ta0)8eX237)5<RcP@5/9&_Ta8?_A+[A=;)96W-J
SY-]M.^L=\L2ffK?ZJeE[>)9G#^cO64Q?OGG[cZd3(3921d1N/S-64EQ_21#E&?D
O8I?-[C)ARG[EEX)QG:T(0PbN1UG?LI/=C:d\a3U_@cDEAEN)\I5bcOY=^gCcVP?
f\?YO_;feI[N#.\.S>#2[I:5:0ELOfGe#DIAF7RGfDOONc5G+O4[T\VHCTH5bSA1
=gN7=Q.._MK>GT#8UA)PdKI12CI)=AI2;;:ET>JeA9#;O4+.d,#ffg69JKPTPMd[
gf#H<31ZD4+L@,&;VJ;8=>]XD]9VU67g).&.a2d.KIWJQR9P7@EBIAQW;IEPT)ee
,&c11bcf,Jd^e9ME(OMgMMe/fNd?)\Pe>Z#<d1LF=e=UC7PLf[S>-+#03c;BI]5:
beI+JBUO#\@1aK0I6\/;4EU?X0&7Y=7H7.@_:;7S;G#DTORZc;&HT(0)=-B(TY/e
,@.4.LX,.7\-6fDR.,;bYa[W\gPO6W-f5;/2FEL-((#M[B^Z\.2<_CH6W]KPbO,\
QOJgOgINJ,_2]B].PF?a]\]Y#f.AZM@07=\CN#/L<V?S^M(E<K)LgB<C#/gGH3I9
e6MR,Hb[&\JP>7Q^&g2OG_CA3\7[1?HaOLKIeFZ+5\&W;db#6H?A6g(M44aENfRa
DL=37,3XLb>DcaG7G5<BF[#LPZI6I(@FFZDFgbRR7Z.1TfUB0^;R?4L>]_WaPPOc
B?=C-A[Z^/RCB@G6;1>[UgTcI&F&:KR0LFZ#1H](>Me3Y+dK_f>c0:<b1VOa@2f;
MOZU23cXG8MBVK3_TOCRZXD;^&3Jg4C>#^E[IU(&TW;M-IRg1PM5<+7=X@:g<J:Z
58]bQU:P^\8ea8UJE]F6ZeLGGI,f/Z=Z;=aM.M]\dSM-2-M,MA&M?#.C9H/>G0&/
&f+A\?dX5D/HCXE&I[).45g6L-6?&AKL8([@;GYDVaUdI@==<+d=6YVE?Y,4]P+8
;gef<d\b..ZBT&OEY5[-c9)T1agdZ<:^^M6:)bLH/\^W4<&fD4IUTOW&(S]Pc9a6
)bZ8R+M>Y[<I0M\WVRI97L29<gCQJeG&6Y,e]:I\FX2:LXGL4^9]cf9)WW\9^9#^
cZHWSf,E2af.HV2P>K=dOC?8IM=0U]^1#e\XOLc&CS?F?YNAC2AXTR@E=:XMX4Q1
JY&NaGZRCb^>=G.PK&]#BCXa>-#b)@bgc15f9a.bFPS/ME8VM7-]X9^\D(0?7TLa
LQ,.V4T(?__aL4J4Y<#;9fcLSDYfcFDC4^a>77dDO]e^/,eM+0&8MIN&FZG9TOKZ
M-@#S[Y6V>JQH;aAX8>V=\NDSAR12=\6^d3+R\Z/DMZZC<^?DL5a1;_WCT><G2L[
YYW;Y5(,@?I;3A3;(V=4b6N3)BAP=BZ9+e52/.ENc&]1L7[.42GYH(L+ZdMA6)LN
VgaD@7ag]3-M]WfTWLHd@;E3=Q>QC#0RR8/\=[X7b3)f[H+eCB[eX8XNG>LV^Y6I
(U#@QTC<8b#V.C:EZ7<7Z)R#/-:>FAc,bHg4bU:dMXOY2RD4VVV^TWE0.FKR12Y=
?Y+8BF&QW0)\G-R&ZON,</Z<ZGM[cM76R&-\RD=#OR+3B;&XMd:0Y9G9L8ED,=?8
&98D.PLfTAc1WM_,FI;7L#K9C^65=30YO5A>)PED,NcFM,HUd[-c@b\gWbH8#B#R
[eRX.-NQ/9E?AfRB_Pdc;YD37M^AF8XR?24ZJ\Q5]T(A7V7,S,]B\HY6TWf6)OII
B+1B/)G0b_YB1aMI9NH(_FcGTLE7dM;eGD3Sa>Z#X.MRCa+F.;Ed#5(J=Z/f\W5O
gFR=ODFM>/WISWDDLMP6gNJVE;)e/Vdg6H-VPa+>-INYVc355<L)S&TCEA\+/B\B
eV\()F^c1a451MaYP>K^U-a4@e0)44Q3\DD61)JU[X21cYF?=^[ePgU0C^NIK9E+
I9\7]8>XD8)D::Sa&]4-\ba;LP/7U[)(60bdeV1fDT9LeVBeZ;,Q-Ffdg^aPS+7&
V#,QE:B)XB+[MO:0:O=114f+KXGMe<&^5P,.AcY3e)#[e]IX5Y/O,aNZ9cGf11IP
<EeRUIC&gWg\[/HP0HS^7H+(.=2,,0V(&4LY5SSGWOB-;@A#R#S]X5#A-/;&2LD3
9\;9V@F_T(@T)B,LU2X,F3@?edI]bSUQP;HfJT:5U\931>?9^PL6Y9R+,S,gbP,W
#SR28NfIP\[<;\D3+OL^LH0c&8P+?4=/aXZ(gTeG(bQWCT,4A:7FaIg:??Jba<^g
VC^Q>d<R;F8CFZKbFeNDb<-D>A>D)ISK(FT&=2#5[VXZF_N&RI2UB\G6^P1\N.(_
T7U.VWb,eWP.J5)QD.Jaeg#;Lg/L@?<E+LGKK7CP3eTGAYXdbDD?DOBXM;552^;4
@?\,R=W9E@Ne9)3@/GYOR_[&S2V?DfaH([B=::505KWC.(Je497-D>AFAF(=2I8M
FB=@<+4f>6[fYDK==,XKUY2_.Xe6\,f==0&P>++6A97(45IA_;f[_=_9@,V-RX>f
A,2EMJ0?64\=\TM\\ZE@g,:CC&W<&B@Gc@(+-30A@df)e.OAR\bOZ[1GJDaF<HEX
5\=Ng/4U8I19_dXe:)>BQQKQ&:NAVKgDd&#WQG#U]4X@MTN0>DBSEb(JG0AK7G+O
UP4XH4<DXL@</8cZ4G+D4Xgb12HS9@&JF;+B4C&:/a@dJW3W6^?D)?A5dG12//0H
J1S=?@HffB;_^5P:UQ0T,P^,92.4D>KNL?D6F>=.N14S,NG./^ab7-TKL1N(PYEO
6a)DPGd9<3\-MCf)TC9^YRNQG/@P<Zg-ZPT3M-\V.bHAcJc@G/4;Ff+<?T1:VO<b
BJ>NU<F@a45.C)0S[W(CLH8QK/TFAc]#dWdcP0(T19>S;4GPRL>.38fF44SFEWL?
7O)O-Zb<;aLNCG?2BS+#0IO/bMVK/W6HCaP;-):9PG#:.YC=_g[\Q6fd0U?]_bF5
8AY(-dEae/Vc0ag2:3eINaM_[C&55S+GNW+_M6;6&af;:TQg,fDGVZ=Sc>>B_@XF
/[.O[JD1[a<HMRJ/88]E?-_A=NIEI]FT,KIbL6&__.78LR\BKcFc6gG;C),.OUeN
K.WAZ?XZ5S5Nf5fYMFdbF>b\<:\T2+cG:TBCY1FH&T.IJ_cR\bg#(-RRHK,<.aRY
EARBJ-(7B2W^g_CQ#\a9]_Q-@Re+VO\dMbB>D]\c4L0R#C4:SQUaH1<LRIB#JP95
WDA0DbTaGSL[,RX>=eWcVHBD^dOAcf.&Q4D_Hf=[@bXf872=3NXZ>MBe5X5Vd;C2
eJ6a]EQ&YD.BW3XMK.FS;52@8RfYNJ(]<>SGF0H:@,bVY]=Bg_^6Y,\)OX?\/GHQ
Y;90[G_HeTdZd96X@.995:Ud_Q7<JU6.XZNDHIU>7QeA.WJ3?+=IPUJFYVVc7[F:
M&bBgg]g:H+_YYc.,#+@_eYb4QJYMTERF_(_E3DOWG\.?)JTMV9dP[2.2T3\_1S&
D;]OAMDEgO4V;>.(&4^OT_R?cU[dUD#0]b=W(@[W=9A:J^L5;b9:>CPd0A,E9W)C
>#dc67EXcX392J-F?6TMR6O[<6ZU,H[7I+#YABA&?@b>Y4Y0HGgWH+S#0EA?#7R6
8HU^6d5M3>OF;Y_F/^/dT80N_1LK)CGQ#G4MG3\6Z;LNdGf@&Y6VIbD(cI@@)Tc:
@+3Ta/IT61egFe7.-#W>:<O[N@eD=+2TI4A3/;f]8M<UNFKM.1YCbLOF3-N4f>H=
:(C>S+5&4XK#:^=[+@bVX&1Q&>_Q?4HO87<2L\_O@U_\G)LKP2d2AE;cYW&X4TL#
\B:RA-SbK&JT_>-^gGe0M^UBC_:\Xa_F\A+Y)>W4(dKW9d)_H.a2_\\BF69LYe^2
)[DG6J0OU+URWPKP=Ca=YaF&ecFRQ2@@^_6LLH3K>cCR3+6-fX=+4\]]3a+8M+6A
2+^]f2G?fFX[F<4E#ZTg67K@OI:;FH^-+&7f3R:ReC:;1?F43I6d&A(B:HV0)V<1
=fZ^U03E_BCTNQ:TZ1.[ZVAM?EMZY5Q+=@2G@]OXO#IE;-AGBWRA-g2D.bCC)\&b
PFfNI+@M5cBAQ>5SA8I==cD0?RYQFCHMXeXV10I61N(OR\&5I<P&c]-R:IDWNBHg
eFPBIg]dO_?4<[F5B,Q7N-WWO,]J#)=fLT((FL6>N&1g@4Q+H:/T=(:TS+(N5VXW
#5IN1>CN\f3@JI_\FAOR+45Ba3Z64@I:OXTa14GG8eg<4&0XNf]QGH6^7YWEIB07
H7VAe:fE\d.0BRM-A1H]aAM6Ad&F&W#F65Kc1+@4]UOP-]@2bO+QD4B):IPWJB/3
aC0U-[bFceEI-b@B)c?Z<&a96@+#E6&N1_D0P^R5?ecd6M&^2&D,&VKMG0MI&\&4
&ZR1Q#XKE?.Y\ASM+^B+(H,0_0GCAVERfH98AVE#@@\SHT;^W0Q_&&BD?R^bY+W_
0gP8W[UT<E<37S9BNN4.)9dKWS1/Z+2;XMLKc#?BKOBK9f0JZPWNc9BF8<5MI:8[
,5>KTDTY/\NTV3/4;H^<XgXgJW28+aK,d[SF-F<AHGFY[_aW;#I.1\a2>2J6SGKB
M8\DFZR2=^YD;@_5ZYZOPb2@3Md4:2IV]CI&U5EAJ(c25eC.F/D#3ENQG9,7E_B6
fM?/A3Y^6#HVDU^fM,g:5^4f:GUfVgQfT6RQZQ)49-IaN0LZ\dd4SQB\W70-?aFH
TG@R]1JWIg<_NP1J_6X5EQML6BFS:L]#-FD5)0KBC4g[H5T=)3Rd+@R9AF4CSJYK
86F#[b/J8C(150^]-AK.c^Yac2(;8BVI@@WTUQb/#eAg.0JC]J5B^dPPYM0T&7ga
c;^_\-29]_2X?,H\)>ZRWf#5a2NFU<egUWfEHg6Q[#4K9=NfXab\C\aL70^IVa=R
OR/<eFYff1[,2\)#U,f#G/<f-C.@W+:gK,UGS=B2adfD)+]QQ]AG(dcDJRcSGY?g
06^3PC=M_T.G4e4JRR)H&=A?](d-.Be3a3g<5I]B68</WH0Rd&,\CFM6ZC?J_>2R
KWQ^VPH8?:@cb@<V9E7&+6d:fS4H^:?K99-B>/^)/(&;5Pa+cSWA_d-S)g.DBURa
Cf^HA7@AL#<#X8L#P+#<6(5+T+@7-G&;=WAUTB<_Y224)gMBF+F3]94WDdJ_?eTX
LL@ISOfO0H8T0:N,#D/:YJ6B(Tc9M5c+@)NGT5g<_H8]9QE/.TSLP+=FK>4-b0.T
VM5K3O4G>FUAV0+SGBGeH4<@SPNV..]Z:#+f(<NV/R<a[ETJ.d5H+I41L/.Q7]=-
SKQY5L]Gc>c9UO\U]@3#)]\9TTC.gbOI)d_&.G41/ASOESJYG2ES/+(O]A=\X1=V
:,Rb\GXXQZJ(LbWcb);V-#Fde[d\2(?/D8aW]LZK);K81->(B:E-#@[/A,.fLN@<
3G/R&d0H&K1GI1&_;N8Q0XIX;K\aW84H/PMPNZ]4VcU45gAD@T1UU3D(=#M+D6eZ
<VHbB)7bV.F/<c6)WJRf_Q@d4LSVKfCV31-AW\5VIAI(.7[/)4V^9?HcCdZ;(c?I
S6eQ),0AeWN#a)PAC?aV9ggFRR+(\2>OfZ[HT&eFe7U]=CeZDc,6]bWJ)^/<\d@P
fIFTX@Y)<g.VP#9LM5\c1\^)c@0<d\,C?(0a)TF+MOV@YX=B8:08#C@b&2)S94b\
73[(5;</57(:&9T,:H,2K6\+,?Rb16(g38DOZ/3aFKP-4S48R_:fXc(()Ve)-VTY
3Y?[&>4^eRY,6QGGNNfgPI)70KKMJNJ]BQ(G)8_dWM7X#,DWfcbd+<A5V\c:;5ZY
/eU62<-^H3\+(0WO@Z?fW3W#B)76:YM&f9QJDBRe^cH-+Y-Y.]2#f:220\=-^A+<
FL,J#bgVe=+c##=TR\(X7V1Y_d2SL.c]Bg)a_\C+T61US2,#V2+Q\\d=0NS:)IbW
JN._0]CEK_5X.@L)c+_>aZ,/IWUGKYK_C1bF7J=\U+bd],[I+STYR:4fX.U71bC0
;_(0#?7AJ1^(D_.HR/S_[9XEO/\10&UE8>R?TG+4E?FBb-g-ba-B1)#5=[,b7_,/
#b2Q<XAS8_J76N(,840JOQCJ6<Vg[L\Y:RH3ggUM(e&C[ED:,.gM)Lg@Z(]JG5[7
6_T=XYN,@fJ6>8f5OgV]cZ\:,c(_KV);(V/-YaOX67)9F(5ZM<H00MgX;+=fe05=
DW=;Ra4U3);B.bVQ=C[#J1;ZT&gXN]7_H2]e;fSKDJ=S-Z./3NQ1OCGfOJ:g->-<
b0VYg-P&378]UJV8]Z=YRT:;Z>O/=;;JZ9)LM<,3KDJ:_N+T4U#Q5?A8D9:BR^VO
@NS\Db#-:M5T_WOR\(40g:aH72E<OcJ5+:V<EbU2CMR^V6+[?A4M[1/[8B9MSfLN
^-IHKVO?PORJG8L9Ie)6HG.)KVR9\F602.6PQYdKe0_[aa)H@a4BY^0@c[N]I_XH
E)cS3<aUW0d4N,F-Of6;YOLb(7,?9X5cDGLWV\7/SHH>>6dcZA^e.-9?,<KNRd]4
@1V:MGOE=AQ4>#MOMI7LaERe+FPD)04Qa@^T)&\M[1[^ec02R1R\e4,#^.b&,Zca
7efdRXZZ(A1;Q2aU;6?P?dC/Q?ZRMDJRH8EVFa>.6_a++ZJeLPg@P_IfR)CL;+c#
GJ?4O9^Ib2bBZJ2]\44S>&eF_V+))B]+1X#<BULA<H.G:UW,M(cIPM9JOe2^9AI/
,=,d@:1RYRH88PPBH/+cN]7Rgb)U.LDZ-V#eU,/4>7,.?P.(=;G\Pb:CN+G,-W?H
9eOSXU@cXMLe/Y5EMI8+A1^#ACS0f\3WXR-#1fNV.V[=E21V&dD7X51<e>eZ8-<A
aMH=2_N2\XQ9Eg[QT&KA,(FS4A<272cD56ffE=2T0H,:4D&^5&0,NLGAQT/VS#1:
PST1#:NUQ:]e2_+S[e)CTKFX<eG@0E^A.ZJ,D477.)]WL4INa&0^c_HG=A&BY?>J
KBLdNBB->eXO5_M4;OB]:X))WIfNS:(_T2UAVZN[eI3,9c449#DJ&(W.TSQ#70Y>
2_FYe,YP_P@]c_V>TZBE7_.&ACCTeM/QgdgaSS\;CFSP</5C)&64a47e77MXfZYe
)eYaT@#?aR(##1)2L-NPgRT74B&JT\R#;+:aT4LD&43MM;7_0aVQfZ0ACEH@A0c-
4KET2<>L)Q.fX(0TNO-G:9+NMZBN:K5>SWc=T7.?<AX,TA/bV:QSBc_F96HF6VP_
,?_2YcV)^>TZd9DO@]KJVKWJH-IO,7(MFTNGEgDKfgN)JE36:TA:S_1GbTBW;NY]
+Y=;a#V@_Zd(L;/35M;DE<#N4E,^S+gVCO0EO9<TB:1O:Kd+8F8[,e-0J@R/;[_I
#KJS&]6[S\+@a093VYNG7Hd3dB]#Q@Gf-(1Fb:DHGO9_V#3@KE98dO,ITR^8d=f6
Daa14^(#UVZc?H3Z5QH@0S\DPH;dLPU1e;g^S_.B4NC@=H)\SVNb&&C8++.9335@
/V_I;gW#L/Y<F7aN4XFG\GEgO,1PfTMPBbD&Ab^fH^X[_bc+/1+?<?\M,a9;FAGD
6C;b^X4P?\]LYKC8A7\HF,#PJDS;G5SMa]BNL09e=1:2GVQT@,7T/^(?<(=]9O/5
,#Ec92;2MINMEag4#1b]YgGTL]P..TQTI0(;Ec[^b.P552<#dC?)Z36UgUZ+G=J.
G/_\15I0(F,#M<;SK>C6-_EWJc+,^[e>H4N)gd6H9O,/.WUF#PQ76M,[fIZPNSHg
9\cK2HJR\HT&]19DKXAgOL),d1Q5#D]Z<(M<,1b@WeNH9f>eO:WJ&A4a>U4RC4<.
V8\0C7B.]&&E-DAZ(6Mg4N2WO[/D:91#&B]?9Z&3Q4^DJ),MGAYAU_.f]-]L1)FV
4]+4:_9LYEcR-9Q.I417/Q##UB>QC[0RJC@MM8V[IOE9.,b14C<3F9bI^K?QS)cQ
BNCL19(-B/8AQbQgI4BEA+?2Y^VBc7Ub..]J]WC\>.Ig=I^HYQ7FH&I-9L965ISJ
/8^5]?Z)0NR=B-KC,YZe,GAc[IVZ+(6e#V[+T_-EA/(/HHJ]Mc15OTJ(e7H=db48
ZR./.7R8/VEGC9VbT?MZ<N4[SQ)NMCHI#WA;V=>==2<LUII)XfUf6H&H&/5JM0+b
K9afM..5_E62B0\DI@LFH@):L;dK6EW\-HE-Y;.OCNe5X,GN58[OKM[J2E4ICSH=
bGIK-g]WfbDQP7NJ+c2JG&P32SGXM&+&EIG^JR59Bd+.R>&10;CW(10P=1T/F98J
2X[I\6VE8Lc^4&,G/#&H.K8IL_C<fPF_KNUTIL0d.f&>C0J:5C?/eHK(A>_SYaN/
&QFMB>GR6QVW\8BG5V-7Q5YZLfWN1?0U+c6O/TN-U]OHG=ECf1C(c;\Hg]U-6@2F
.U,[ceVUJW54;J_@,14)8aId2g@<+.b8H.6&4<W5J,FWaS/9@&Pg0JG,-/T)B#F]
R>LH(e0B9bB9dLNS)CFUZ.BN?RVcC=&R5W;aNRG/fD#Y>dY4##C-gYI1GU9X8-V@
I6O5.ZfK,L_LUB?bDJ,MYe#geaBSe1GTV\+U;,>Pf[a36XPYQP:#5B(2BZP8\]ZU
<+A=/)d<.Q1;5cR8&?-)db/_4#ZEaRa0R87J+FJHT?HZ.62G9VT67N6QTIGE[/T2
,)OY(BIQEJG[7Se4]#SU@7TM-dL5EYJCL<bP8U1620E\BY:U_,_UMEJT01+XKHI>
]GDdPR[:4/+L-JR.)>+=cR3CRLAW+_F>..ZUMFPOWN-REBBQ(E2e\.8b:d.-f[>B
fdXJB0>818Sa1>5\7J]PC+#3K.B=OecX0Off&[#Hf)A?3g=XcHMNTVQMNfP@R.g<
9-SI0.L#,GHVL[ZML,ORe.;394S+g.g^IX1MR:aJP.HUdeJ.g,U3GOW);H:O<J8G
6H94I5BgB895g,:)6N-GT&#(@U194_9NUD,Xa?:[_-]Gd:R+RGaV_N+_3Z[<8>bK
(RaA(WI,.T.F5ZE96;+APN8-C>@HHa/Y12N_)7O,[@5<<DPIORICEA0PeE02PQ]Y
^/A2bg<Ae>/V8X;43ZT\M&FE46E?0XQfPA8]f(a6PIfCP&BK_JSUB@=K0bge;&;?
4,X+ed30Zf#VPM3_DIV56f7d]5#2;bC;OPUaC0)QDHfD,0;96RII,]&b(#C/M;H7
I7gT8^c1cWIO[1;S&3g?II<=8-#_b,e8/F+cbB5>EgB^9(N0[Mg_:EU0+ZQFeX+N
,_=N6P=MfCC,=?7^7RA8C&47eFg;U#;[KTH036)cAQ<dS?Y4>Ff)&)c2/=1\=)[+
Y;(G>-R0J#<2Z&VR./R8\K_7[S/O2HgL,N5U9C1GR?XP(]B0.QU86a[6g>7.;DGO
TJG93b3LdK@O[f+(G[JQ2a\TJ=#3Q,@_N1.9P0++Z^J@3Sc<M733Pf,SZ1ZWC@+<
E5OHDcGIXT?,P.ED-#H3[B]fG?/GTK4)X>3G_J&.-B\g64YQ#]^D97PIXcNcY25_
BQX9Y>ZNHTA,NDKF28Q2N7ZR6SGDY+R-6bQ#ZHU51JKcD,N;NOTa91T\V]@T,e8N
.4[;4E9Ya.e3PZS?33D_6GF?I6G(M_^A[=Aae>>66L]:d(_4Z2.=0:^f+AE8-1]>
=^8Zd#E]\QJNdU7WJIC^0U-OS35WW;482WR=^[P==XBR]);DbII+-PT)7/F>E<c>
SRW);D4F:[55SeIO()[H5M(.@]VO<GW=Q1S5YD[Y3gEIHH/1;YHBQOMSVZNW+M@&
4:0>P6K;IQ=XU,37f@2\cQ8DFUbRSX.@eOE:=5G;J>HV2R3XQ27A]TRAWBUPS2Ra
[#0SZT<[(=M,U@WDY2L+7+(a/6\IC\d.3U34KAAXHA-Q?M8#^:X0#F#JG&HVfZX.
>2ABOV73+I352NWB(^S3EFC17C<Z27@61@8#QL@=c6TBW#M:<:g&L6X#a,L/<IS8
--R<Ga--&d#R2SX=(A9dP1#P[3,1CLV<OMWARXB;&(Y&:_@5K]ON./TecA9A,<aM
1UUbaJF0@ZK=LQ^&@])7f5Q-VU<VAa2ZMN4#aRE33#_Z9BIG7^^[fL(;I2W3B;5>
a\XMa:(a[b^@6EUQQf@-\Ja22#-NU#Ee/]QdP,&V42+4[N;N2FYRAcP5R[dSaL_b
W&JJSR8:^YSM[>^UGYGF2@Se@c]O7SZFeVJ1/91SS>d<+4_aZ)NJOPL-<5#b3(bZ
&Zb^>GYSKTVH.#^f/J\FWV_IcBe#_U\g6JE/Ye4;3<bSKPWgXQZYXbQO]#DOGD9=
eV+U7:4VSA-a;.WAcG,WHa<)adKdfU,cHA2dRI+OH9M:/P;fPC/T;cDGTgV:\SPg
+F.:L\3SMBN9FM2R2.[^#B((_(I/c9SbLMA&H2/[+bIL\Xb7<BM4gZ;70dKVf-d?
?I(H&HCc5>-P5QB+E,@36T0UAbWH;KKaR2C.aYaP=EU,H<cf6S<1Wd\C3V)(P_/1
OgGBG_Ab2Q=GFY7RF4[,JCJZ;.Rd@ReEJPaI.U=_I5_8H3a+QScM_g?&=bR\\A#W
B0J<^#>/3-B09d?.ZFSF?:gG3(@aaD5]]fF?VIT3AETB9AJ192))B6M)5(:B>G.N
AP1R?,Q-VW.P26.a52APX[J7SbLEgS69cW\@\_,Z()<GP9^Q584BY.IPKG6R]P/[
^d)S/R8,\gCZYK90[7gS-7A-cWbTXH(C,2;<6Y3?Sd-;C-4-XLZ/,#^-RPL?54(H
b<YUSPY08^9M-fD2OF&d4?V9N(6<TZYb7D41Q+-PHD;2VS)<<eWYfUgGY2PFB0c/
>1X1[R:1H:bKOgP4;K_b@6aH<?F8B]a(DS4_LLYROL?F]=c298N)#gC(Q3f3.J0;
6cETK7^)&L-[C9W@;+).Me5ZZT(d4>/CMNI>_6@:4A(U)RVRgd&fWdIg9F#:D(d4
WAT@D>VX62VcD6ODQ,e5<OI8MHYI)\X(fF1X-P[KXC0&SN3I3&F(#EV[4ca0K+2#
;M_EHW)R,E&.6TWRYO_1af9:N_P^M)])GbDA1C/?SGWR>/fZcAdac4:fgUV]<>?5
N0RT.B1_1?]C9D:MN4OV&5eP=Kc8CNKZWM@?/.Zc6]g@25EII5V=_+CBS1+BeF)@
4;ORFDSRJDPT)\I5U;/Vec:9N,d;U6E9STg#6g&bEFaUPDBIKZ1R5MUD1URf^Rb7
0[WR(NPUe&HV0BRGa,]U?XQ:-4&7F<(2FCO_KHdQN.=O,5?4geH]-cSD)DO<WX2L
<KfdT5gHfg5B9Vd:/V5/>?J/;9XRJIGN\_dKV@@F>;27)JB,JZScQ^FJ/Q\?V(Q9
N/V;DJC-+C6&X4_XD/V>&1d(G71;WNI>;(8VW#[YH(cW]MJ,A+J+<-c=N:XMW?cc
I[^<a1>dH:FTU14C[I0[.7+Q;-fdMc3K8&DVTRHb]607((IW^\Z\YIN4).TQbSbC
D^G,2W-+1G+_?,.(3df1=M1U(&F]G@eV<d\6;0ML5DJ@#3,V<84STH)VV<<>(WBZ
g6G<CZCec]&#3U#CdNf;)^[a0N.41B7PNYgSZdU\UA@d]ZWA#\T]-)d/H,6F+P_C
86-bB7e.QQ(6&VW4R@WX2)aEQbHK)(DC4b_W2EK\,=L.M_RYW(FI&\0Q2N?5#41C
&TQ8I0>=SZ#QE\(9>VD+\#PH=OQR]?[:5,S3XP1d7(<Y/2?0O?e,MW(:)E1A4;dO
S/)S9URXTb&C]2X3<d?&bVN;2^X4877-DJ9&+MRX&EgXBD9=>C)[O_5318ea93WY
L(3efbD(#?FHVN=bOe;<4PF9a7.]:+@BS(Bb+e^b;2MC=U:gSaITC0a#3FggP;eJ
_(YW?(4NOQHC1;)dL<X,+4Pf;(##M69EO>719Vd4)LJT>A5?,I:Qa[MGWI_T;SKP
7,b62T->@99a@efHc/)d/PU57.fT&]B7<6b]A[DMV8_=cE;#=G]?^6BHD1;/[;SK
(F93K,9IfLRTPES/C5D:TNB<IDN9a+^E5aS3L>H0U@cI24F2:/M90??3-c<<V(>L
1BW(,2,d;g==ef>:cQb;>/DUTEUB\X+9b9@7=8AE7e-S)0U&_P8I4RQLNZPGBQ84
W&VCI-,K^>DH1N^bZ<GT>V<ALZGgPb413=]S[<J2HA4[cOM@FZT-eX>9fgV3FedM
G[HBZGNO9VbNG4X@(KJJDee/a_.C)_^8+ID..=&7f,aS;UHS>8BZN[-8-]#.45cI
dE4#9-K8Y^_I>,F2-:?(D&J@Y#N^A5g61VB2bEcG?;8F@SF&F0?,79&gP-g_^_2g
Y4fJ9DW5e@aNI>LQeaId,P:#.ba\?+]Ra;LR=6;2f1LFK=O##g]&e9)XL6^\eAY1
7QM?T2JDD+:NIRdR8J],dcY=D(N_9;VZN/RXF00TSc&G;F-4(?U^:7/IJ48HgK)<
TU]V6Cd@2=Q]]2;B4Z2SZZ3VTVXK@K3MHSe\aG9Z>;aC5^+5B&WJ4K7(0^O=S[[2
aKU,,/KRA&\MP+B]1Wgc8)O2Ec&<\+R=B+c:7Z=S<f[LObGXOUR,(Kb,_(O-0)BV
_YW;8D@\Q?,GA&M(SV<ba\EXRX>LAI\EQ,+HFPaI4=.BHX0YRABaZQ+MQ)Q6d]/S
^Qd?9OHRTN6daI#G]1,-8B1+ZJ#EC-[=MJ]>6LYbT7U.Y_,Gb&JR==M<9GY:/@3e
^g#/-6^#(#g?<fGER?c-24g9@+G,>Q3/G8R)bb11f?594@3</BK^EaVA3?95E?K5
&#QZ.9XgHM]-=JVJgfSfMea+NZUUDM/24>RfR;:CdTGDX@PQHRZYN<K<256O,<NI
L/N.[0R9CLR+c=fJA0J2SBAO8=.Sd=F@,FSJ@RZd>&6Dg[@8#.O+=b6I7YOQc2DG
.U/7NN[eYfeg&MHCCcOgU&&K16[^I.RV_Y2<17\HPcXed8JMb?QP<7bBe-&=Y9--
cXe:9]Vf[,85CeJJRaF5=)0Cc]]5MMTIdWE0^a=^UfQ#g1KNGAO4\gOCE<&-,9>T
F)XF5)eIJNEQ>JH5NMf0?UY1d)7Q0g8]QR?MT21bH/,<gB[A;(NGR_gR6G@OT7Hf
gK^X8aLf7[Gb2b2B^ALYEPA_)^RW/eUDV6A6EDPe\egd.Y<^)U69UaV([8V2d6YR
BAH=4Q[bdOQLV6a#aWB(QB:I[6^<DI8XCb,X8-f#4K9=PA<E\ab6MI8[2K+Nee8Y
W]UCK(a33@bT6PB1OfH#gPQA>Zg0&<B.8LM^<V).CE-E&d^<W4Ig-O#cMgf+<?Ff
R_25&M0[/V@?WVDd0H>e.La5?L,OQEE&E]d6(4_D<5XJF^L(^6]QB1+1DSKTI1<@
14,(-Se1[]fV^UV>e5I56WHOX3;MJ.W]\GC)NbgHCX+JaMX0QA@\3_e>AGEBb?H_
\OgB?AR?XCKGBM^M@VB;BSBO;fZ,?^3J@J;.8Y]DaM+1U.8P^SQE1ASH;G:Jc:Jg
c.=+CYL8^;N#6RXQ_CJ53beaIWaN@Ub+19M&N947,_+>M][7Y\#2.gPNM,2W#dJR
ALZ)bbC]OG[7=GZA&HeZ-4=@<)3,-0H-R0^(=6R5]g5:Q8Y&OKD\UBJJ3e@(CWeV
27JbgBRO7)I?0WF3XGRT&R-+;BH]G;_CI>X?R6d.0)C;.deL:4>.+[W3H2Y4\;a/
#M0L<ZR1f])O6BH;a+ZdeIO2[>+S(;JKM6+#6SX#C_\.E_gfVf.E6E#N0cAOFN:O
G.,VX\7GJBML?0eR<fFY6]AAHU@YI4F.4.7,,]IPeH:OBPd-YO<bB]TC>9#14;PR
D1g2:E&7CK_WMJVXCEZ,5.7\,9E@^NB&@4(40e=AdR.PIeJ+K6Pg6V@GJcX5[TNO
>0^&:Y776SMd_Rf-1.FOB,1]PCJH=)6[WQ2Q=3>R&V^M-N8a:4+>^A\XA?H=H,d3
@O\b[TA:@WgE+=@/QF>DKVcL3.X^>0)HS1b3-HZ)L7Y_B;^\CAOK=&)a;9+decZX
f?fBBP;-FDE.]H;N=4-G-g6ME,<DV;aE^BKe#K@D<>Rf89;&_?8AIW5M7BM6D7B1
N<))b696YS&&L6MgB_R[ZOL;XH[LS)?KOCU-9C>W3bP2CcC=4V&+VZM.&6,a(JX+
bN?;RNQX[^QEE-7BHDXJD#eQFHXg+:]MQJF@J-d8DCR(QcZ..V^M6T?9.T49YZ)/
&EP49\#IJ3GZC.EG1GB+)PLT5UgC)X1WWXcTT6^9Dd7T2F;P+Ea_I6P11/S5Q\Pc
O?H&5B7L7]_QM(-TNd=7Va;QE+^=;X<]C,]C_URD\4dQdPO#-[2L;b4=X#>(@.OP
BU651^+]TDO(_WO7O9cW:.=14#[9D4g2M>c)[4><07[5N#LEUd6O7238(3E::<>8
@)\79D<0E\RX>\H=]R+CKd<@ZEK,D]U/V5H3.<;cWZ>OcI4e;ML9#<IeTZIL/^Q+
ON?Ae9./WX0Xf\<(8C&NLI7W+9YONZ#[TL<<P6/gJC2A1JW<cKQC8g^Xc[KQOd1R
;85=.]32I@8&cge7L4+f3@WNYg]?9b?)6PNVN-]@?BE9<D6c6A2#T)BJALSdHQ&8
-gCTCFUDaCBSeC?&e7/J(L76ACLS1L-#_ZPVXFeFXV0Me^?0IH2V3ND7K6UO]K]Z
H3e.?Y=)IVSgXb.;7WUF;<X:L+8XL>=X=GNE0/DEXVC0c8GKTfM[GI=Se\a=ST?X
EfIFbMO\0Y\1/47AZ:&N(I=M&,F/@?X.JMMYA\g0<N<IOUfbKgA7/e.PCgJPJbHM
L_eZT]P+1BRFOaN@VBE.YRZQ#GWO)C.Q329IaE;@IDAa5&C\L=74N+KC/b?[>.C?
+8X5@XT1HgMHKBES?5bAF7:ZGe+)Y+@;VcSaf6YWK_,gb?c.DOg.Q1IY2=^TN@OX
(\dUge58M4#CA=9]49f-#Q,;J;->PX[\/\#]3(0/7C<END;[6M#K;2<2K?Ob_SW<
--Dd<MON-IcFM(A:9JM^?9Z8a.J,&XS0b6,gF.UgH5:A@[ENUWCNY(?@(]>W/&H\
._YX)F#I:B?GWC_S/b6ISJT5Kb.\eW)aJ39OZ2Zf<c>AF)PV+eWf+G7G4K>6YYWP
].6bE18Y=f3CY_),LG@?bKUX?UP9LD,]dBFaFH?Cc010Q@(fSMF9AU=MGQB]<I((
55^bVRITCT)M9AO9@]3O2K&2A^?[9QbY@U.9/70^Q(74P6G:8^<H@P/74Y]=6.&M
=W#4LfT;32N\WEWe7I0?[MF>ZZ>P<0QQ4D9>]bBFH5Hc>f71E-T5)=-;&+5BX[#M
D,L@19?0DIaXWEgE99AA#2OP(ETa;gW3XR0T)+f@Rf<N;DaZ4dGVB=5aA5XMLG^Q
S?Q\g8Y<a1a]b>4g9&J#c_bJ3F7Z)P68TTGW_E50I:7I:P?fA6@5H;[?Nb.)N<G#
&U]@1]_9]<+[=FN+#)c]J\Y0Z4.<;PV4#>bc^@C2adIZQ<bADMKBEX@L)9L;aF@(
^UT#Y@Qg&@<.-e:TNQ=+)XDI1&/6\aVcOb,5[V\>SUd9#QbcJ:Z.\79Q776/._E4
TW^CK=5JPKZNdWP)1OYDFg2B(D<GLAIXEaG[/COW0efHC\IO/^IUAC1#6=<a<@SK
2YJFY@C\:<1L/P?0><2;O:>c.WB>Ke-c+;4?P(+L[LD7?A2Z3cRE>_NdZ3-R]?9Z
M-cLDIG[:XC_<BD6@dDM/dD]]3X,KKER1HP>^Gf#T3=<PQfRFUAJ.?ISaQ_3<.6Z
B??FWO;,TN32]5FU7.FKG-aTYY6R.JC+,gAK=e(e]>a8,c#&[A2EF0=a#5=D]1g9
IW>@DNa59172ET.=,8QM;g2>P&4]Y1V=/+:]J@S/ESL=7bJE7bSQ)^8=A<@EJBJ\
.-KRVIU.^7GK]g8&VQ,,4V+M8<-Z[@\/>d\EVJICH&eX+>O=>1XK3fC?IDCHP55=
Y52IIEM52.L;58OWa.Q6e1JTGT^(Ie.KcVCgDFQGHO&;LT&3ddeX5NfL6[4LOV\(
0Z@=fS5Q3AS;F7U@4+bQ,E8#ZNXG]Y2VPd41)(=K#CgDX3PL_8E;;^La]HKcIed3
#=RB6L_IM4<F878\c5\c.&3:gC/WLbg6T?0dEg,[6MdL@:J@^Zg-<JFI7e)#DS5f
34^O#_HD<GS#a3a0dJ;Zb:NRc@Q>f;=6<e;/dM;bIN_LDEAZL9KF0=fF7U0N5YbN
49\V@Z.=\cWcV./:87V>FJg_-A9W/9.B?()[f89)3/.ML:K+6I(V8I19HG?XKe9O
ZM2^#EFV5SNgHK8CGTC5G:dDIM5;(I8PX-AAD:\W?bfg=^?a_07?_3W?^[&d8cT^
,:B1gMg^>\Ua4P](fVf<b^c>LU3?ddF/)K2(LOH,V#CK.Y5d<&I1@d=-\bXDWU(f
;>-27A^1:LcaeKO(:-K-2;-gXaI4_6.Qd+/S1@(Ag,16Lf6;T.]AB.J,3A8JE\LR
++6W=+7?A\C2[>1;=-DI17eSXf6/VGUH>5,QR-]>D]W+9TRfe00CNNY^f_+g15_5
.4<4ETS.VgbR;CFH,2?ac;G2<F]7YY/7H;IeAOd_(ecLbV0XgT+1<8P(+Kf<b:.C
^;0a]/L#E;)fb^@+\&AQPQ9DJI:KO&IHYM)LXG^BHN9M0EDRK3W[P2ZDE^\AV(94
]\R-R[eVO-gZ7C7L4<,RP7S;[]SNeUP7:94ZO[.]C3.,>\O:>2;Q2.dU^W4a<[PO
d[H,H>R1K@R4<&59>^](RC1N[O)/b6f0&S?[PGH(\>;[1GBcNLT5RS,W>9\ILMW6
:EGD3Qa@b@:5[XF@TS./MGFS[dR2IO#Bg[Y&&Bg<cJK<?)Jc7+g?&P;FKNgeC;<g
EP<T5a482/Ed>fZ/.EL(F<K8TXZ:/3R5(#9M@NJd,b2+O3\L;D26P;1eMCB02bH/
KO]Qf.eCdYegF6YQ(0-4,fgZ#O@QE8f--WJ(FIH]:@B0Tb\CWH2V_CWTBRcTJgP[
W-36XOJeg56RP?)b]DN^STPc^fVZ++6\eEWJ/PH==JN72<K36?U3V_[KV6>+(2]Y
a=MS=<cTNOTA(+QI3+VE-6B@IN@XAG=>gC(71Z:.R2;ga/cUXADW-#]J5LI_-GO_
9/Z:F]_]9)fJ9fV3Z>bLJ-4O;6;__<)8H,O@1ZT>&IUPb0f#52XBPMb+ANX>K?RD
NN/M.DRT-C,-M+a;QGdF?b+>Z4&dX57gN29/(762L5,5.Ye4#gTe-RDFU23PC3B=
OQF+5gUL,a:g]S2-/S:CVA<7K12Rf)D@ZKdP0:df5\9d79(#EWFC4g?UAHgPS=f5
<L-0,6?Ja1Mf+6S,\DYP;&R>W6YVAS5@2>CdAIC&e?8@DP1&:UH[Ff)KH0DT,c?D
+eK&eS44VTd,Q;a.]1UT_@g/6\VMd7>b91DT?dV3b6#T\e?4T.D8G<9dH1SZXe,W
L-R0/>aAEMdQ2>+0,H3SZU6,_BHgSX[e[LAaQ@?CeeU<8(J(X8=2@1+73b)QZ]:.
07B9)F]66YT#,FBE+>f<1?c^-?(a=S(X^]^QMfT:)+1WMY39&UDY8F1/bT,;36?T
W>)O&@O2?.M8A3)gG_JK_-4=)]]=V8:;Be\V2J0[<Q82?7@g5]DGb85/S=;GUNgI
ISN#.f^03<&OgXNBJXWdLU]:VB0[LWae+H7<c[]QF(c7[N4fV\HVRdZPAZ]O=K8Y
(0+KID21_W_8@d,V@@((P?6)=LQ2a0EgB1=aG+,YZKYggEa.O3)a1)Ea>:4DRTMD
M7Y=)]Y3)dgOf4:O@U\&I(>?b>b\VSU<EFVaf7,.bF]>c)Sc8;dYegBM9^KES\9c
Y3\XJ\,fJaF[S/gS#FEgc.SPTB<0#^\7WI?a7G5CaW;=W^=&&2KY0[DMXX/V[7I/
BKX)S:(gWLYL;>,96AC.2JLJ5&P::.^]_BMe;IX(07e=,]OeNd]I:..@Ed@GCX,S
Ug8@bKRJ,-V+e>/Q_<WE3Bd^H-J?dSUdSb0_U[Z>a-HDb+K#O[Y&;3W#M,1BBUKD
AAIHMMf?W(,c=]-JdP2S2:,Q>/+<)f0+G/[A]S7P;C\Z(BKH7^KL]aFgTB)JOUA9
^Hg:aa5/ZW+aIOHIBc\cC)?DIecL>HI.b\g3GX<^Xd<NG&<4HRG=//>77&2X+OG.
-9B-5@UgDWKB\.d7F2QO/MaP&AW;fFFNg4U\#B,bXaAJIcLH<#O8EK=T;--cFbfN
F_LB9geN9;:NEOC<?^,Wf)K[>5:Z^WDU6BSQQS_7(X/=;)7ZI53cNM8YM91D=0N+
E:NO42TRXIU3N0c[-IQfWR^N/.KGC#E5NE;b50XfI.+NId:\<CbXJ);;\aPG>_]@
;B9efOW/@QgA?cDQ.?(YN:;5>d+QS/S9PUB]A+eT-7^1(N-b_PV]3I>Bd\:fV<K[
<[R7H]d<YY^F?MG.e7RR]_gMN9(2[YYSNT43NMV/PKB:(87,UW>+aU5ZP>7acRM+
UaOB6O:QdcJ_0cK>D7^S#c=-QWS\+N<Vc+2#2>(eRIc&5>./Ld._V#,(M^&TdHVL
&PQ>[L]RA<]A0UPc<W[b8/)c7VCV8N@@Y53U3W9R]HULd=F6#XcOc/-a:/?HZPR<
H(a4Y#UXJf1EF3ZBOI:71NV3#_Y6NEF?ELIO>OPA/TA88Ca&HTN,f=DNgQG9W\YT
d9ZdJBOB<D:1_E7,gB2<8dWTR[5BC5^2#,_d;NZf/QLT,b-)RU7:AcCa@F-g2JM&
ZRg;#]LD3<\P>Z#Z&=-HEUAa[3Q0.6(2<_Ef@K+e^[b=N/POB4)bF11A<d7_,^H?
@Y^aKD8V/bRYAQ9=JM=0XADKZTG>24e]3Rd^7f<DJ[K/8L,_3NDPCA)Gf2J1+1.E
X3/d+>(Ca&e?1MgGH:X0EO-eZ3V7+1>;67WFAS)S4ef71>V<F+U6N^])cad?V7Sd
a]S(Q_KWQEW+\f\S.8&<SaFbfgM.\Y0b=WWZbT6Z?P^R,SXBf]6^_BgK24g1F=R@
g6&++Y6DO,M_\D.C9.FA_SP:af]3N?OO5FM[fU_](J.IRKdW5C;[@32UKee\O0O9
4J\?aZ3gTN:Q?,O9d@JBa_bF.^>?+9WF4<2Wb9.f(M:]fE<(1IKSGWA^Pb,#1fJD
CUJD>>,L.3P+3Ibd0&Ig-Y6ZVOR-B6+WBRMY/(@C@T,.D=6A[aO<=E]/;7:R[8QK
Y5;NDeVYOF#<VV<S?NQB#,^W&_eSUCe6e<CQF[bfQd-e6+95BFB7RR8W=@5FO)52
=ND\bT<O,;c5DNX_0K&2^bUFccDbFIaHND::HEB.0KE4]g,Zec7cW@SeDM6d:Y&;
#f@[?E;gRBFTCSaVeKB[^F#dF9ZY+aQ2+J3I76OS86RKN3BY8(F5AQ0KEP@3VVbK
EUJ8b/HAa4@(Z&&?QEK2;K;[BX[bfV:eNF90HQB#TXT\788=E)LZ1BeJSYQ+[FB+
GbP>PMX>9)VLfC;3:/,/FNM-=<K+-9RACe..9)BGP:98H1:W:=bXBR^Z0(eKH&B<
?\]Q.IS@A\^[C,L;#J:\HgMZUb6RcFTQ_QV>ZTdLOR(Z.))K4_S=Yb6M:XUTIPYX
GVcV+a8YEB6QWXd^Y6\<6E@FLA\8^;GI?J0LUD)Z:<#N-UAWFbEJb&d?(XP+e7<F
F(]A)QHPD:.L?912(PQIadJ]2DP&04.Nf+d,AaB5FVF,(e@WP=c>V[81bI2-^8a\
S^#A+6P\-WQ>M=GTd6E3L@DRNX&cF=Yg?3T4A888XU&(D-P6#Q+2a-H2fXR\2?CL
D@Z3I(ZCVUQFT0<J5+J(8C(Ga/dc41FQ#:;9I[+FI:.52)_67,+fVVN^^(4&fS8E
NU/9_&J:5/<Eag,f2+.Ca(,e^ERC9CVL\;a3NLcM+6A?0f3.3eb>OIg0Adc^?-@#
I)a@a,65B4a;[1fA9=fWZ[1b@C,I/HM=[I6R?FKTc@C@GD,NY\O(C;Y\97cJYe[Z
_73?VIJ76JO&@/:+O+JGC@_>P[d7P<>g(^+bYH:#32NTJ@H2#8fHM68-,ffb9Z8+
I1d?:_AK^8QcE5c3a3?SDaf0&0_/H]^F6U71H0\MWGfUSYXe)T>JNIP+:gF-NZH8
Z:373]-=8.(?:1d7MY6(7_Z2bZJHeNQF;Hg_4Mf10I,\+-g>BJQKgU>bSBHe\/7H
dSCS:Fa4;7C/H>@Z\?^2KX>>&A-_S-)B+=OaX)U:gRgY8Q#(g@Rf3cA>T1.-@.B.
>F)X,K^1SNQL;d[3]OF@_A&=&8N:VXH2dECYeC++L+(4V6?MP20:+K^/S/9UUMV&
b[.=LVYe\He,/>-YZ^g&A?+1L(CgaX[()>48P]=.W+_3?T7+TLS1QC<XA(S5LZD<
34.Id1\4NFV=)R#3U/9cNW4e?]4QN)b=Z2g:=U6\[YM77>V3N#?9C?CKd&RERBAf
F_RHaa;6O^7>EQQ9@Y=\[UWLee<>NNf>=^8Qed7G&YKEd2UYW@bZ6+(2(=)U7,74
@U?VA+JHE,]e_C7U8Nd]];4:2F?TA3PG;H-bEG:61Lda\+;GfKV(MB:c^dPUBHGP
ADM=>d7/,Q018H91TcS=?#=U\L,-S^>d2:/,BU/cMZ2/\_?9>0WYJ=5;C]3L2[Q0
Hc2UUI^a+#E;dJ()3g<.,EfPBSHKJc4dGONP//TP4HW<2KP?<AB>Qec#gPgR)ef0
>W0(^[7b02&QQ9B5+1<d[d.<&f^W/P,W&VT6_)MR2QdTO8=,2/M2GYA[1M1LEG=I
6WK^[GC&JJ(dULTJb\DfZYXJB#ND+LM/_e\3IU?X).<gRXJJP.V>EEMIgJ6R/C>M
5#+b?[0.C:H(CTISQ)VQ:@#)),<[2I):(I3OYS&H+7.=IHAU>Te;3WS&eFT23,]V
fa@V&S5&9^_/[M5fI&DA;,SED9]PE&=G=5234>KG-dIT6?8\EX:Obf,2<7TF;IaI
QO)5EU86^,2?1bcY0bOA]B7\J(d64CU&U0>_(5<A?#/(.775R>-QaX<O[I;8\LHI
K+:3TBU0(8#G:^G,b\<Se&16\R[dVa(_()_4#-afNa<.^^T3aDR[7S2MN4XSM;MJ
Ncd(D)f?8?-RU#HRA38We@_PI-LQfN(>-HE+F#V(R-.^e5/YLT2g98ZGFdGb[OUc
IBYDEXg@.Ee9^ZBIV_09P>W=3K<O,;-=YUY9?Ua85cO6.Cf.KPQ^3.U)dIWDAO>b
#RO(O-;ea9@^(F3e_SXBB>]UD/Q(.NDRGf^TbCW@JEDP9FgJWa2\c#b^=M2/BC-6
S>Ma;;Y;SCb1UOLE>YIR12KFDZ[+BAJG4bb=;B(9)?_Q^<5I?KaI3ZTL_(;XE@bL
;@S=eE3eF8BLY-I\Q-N8_.?\7#);K6?A(&8F?8<HDKDc;>BS/VIO0Z;U_N6eOf6<
S,TK?;+-D8KEQ.OB.Tf@S.g:fOTXJ4#_6U7d)Bc;FeA?a9:d\a?Ed]I[[+P:E8V,
R;[EU\PbN2NXUP;S[3IMTA+KO4?BS@.Q=X;V68JX5KT+,4Gc/>:ZdXOUF^Y-62+I
SM,(RG+C=SDNBIV]=UY+fg\7aFB0d>IO;KMgY?#W<?B.Te^FTc7M&WE=[W5dI\gL
OSWfC2V&[N?_P);VH&b]S+.cYVZT+Oc(fMEDYLM_2Db;ZX3S4YPNO-)^T.6H?cNY
&X37QWGAM,P)Q6fa6A=fY4]N5eM3PBI?4&2JNFZ=8?.+:K?YQ:g]\@aZ98g1?dg6
T8F]<gVOXcQD<AT(2D,efOP5=?[=JPX@NP;LQ[YLf-XQ-8KSLa^aA2[_GVL#e7<a
QPeQSFA^@a]C4ZA=1>PE#<Tb6]#(Z;K5R2&g-5A,8;-M)0KP.O?1-5-ad],@RMHZ
IMSWO.Z)88@A>?VY3VYGON2XHQ,6,UG\SfeH(-Y.Z=KYeW^7Te/1FYcE96Ae-D00
?G+UOXJS/,MDGRM01RK/2:-)_eIbffBX3?>&J>)4Ba]/8WQ&eW3^)9_[2BMU9Ig_
b;3-W)>B(Y.RQ^&a7_(SX9S6M#4GFOTG6]?eR-SH>-a1D]7.XW;@FeTGOG6K7(eG
SD]/,,87GN3CJD:3Z<>G?]EdgH9ge<;V/RVG:B,1-.MRC5[@;WSf=1Dc]]-g_;f+
+)LR[Jf=.3fFMQFQE.\eIdAXD4.9_)[#aY-BGRAbD2?695^5>INb5)K43YSa@K@U
:YGRD5KILWGH/PER#\f[OZ=D^_/@#_=\_Od3X\BcGN491XDL_HRb9RC15#S(+RG.
WD;ZR[S#0f2G4MNSS1aRVK0N].#ZE1;GX&_60/PI:T:N_>?#-8B092KXd]bF_:I3
UGcKG]T_+V.5,QaL8HWa@3]KLF0\5H3RIS=:HaFKJ?a)6B\X+8d\EL0SKdT\7WR>
<YASO1;d2^,=;W?[,egTAXN6dW(TR]\[W.])/ZR;K2N<V@3gY=\Gd<S0;G9c3+[d
8DS8eL#MIW3.F.&S6?+eD3(7-f^[?LGYU-PXFH)Q70X&J)B-1;_U0S:=X9QM^cBN
+aTGgI8W?FL0&N3W8dfF7TU2]A?U#+<@E+))bU>_@,J:I)]Xd\75E_,^:^Z^3Q,Y
(Z=SCGHEX>NBMH?LL[CI&QG>K.V+<DCS]]f<A,cc:f,4ZZbPUA4KEY,gUd#gD;>X
98^,1=:._Igbc/f8+B5#aE<;F,N,B4&9\Z77ZD8BT<6gV7;f&EcBc2LQ0ZTdZfZH
19W15Ja_Q)\F?RN6;M3JFe+_X@+K^R?OYO/Ue4AP(,cI8X9=KU5<-G)>Cb9SIG^2
R>D.6N1ReW7Q>K2WIL^,;-UIG/3I&3c\^<;[)5BZYE&\fRI+&=&VF0KTEBbNIAD#
K1,E]]KNSQF8M<a7M#/36XLYHOdR>+\@PP6D[UB/R;7RNf&^+^<4SL.B=02[2MIR
77<4>TNY)C&[08Na@7S2RO86VcS7c2;e[^]&[BXO#HN4(08c2X:O#S;+:+@QC8\6
?C\.F8?9.4;JC+JbO=IA?DEQfSI<gDG#\]GBE/7TdO=K6A<8WHYLI07E_.cVUBe^
WeX^W.Af33DRZZ_/#;1&4FP_(JUc+(;]V4=VMLd+SS\O/cF2g(1g4YNbLOL:R\4D
<JQKZPHHG?;@F4;;JMV@Z\BQ(@3ZM]XaYB19493d=AIKN?VXf>PfS@+J=+.:A6)b
R>RPbKX>Y4f?E(G#]UcUV;ZKbW3/_6H0<0b_RLIKN#-@WK3H68\b?c\.PUEZ?(_C
-XL82.2Ze1MDG,(G+BO0N.R.JGS;NK7AB4F8P5-YOW0/5([c,?IUSBR38Y#Y1QFS
..[7I9:FR5UF#f7Y?)1-:7C6,9XO(L0g1<<J2S?VYC.:H[g7DFPN.EXIGJIK_6:,
G6I-2KV;XIA(dd4fY1G;J>\DB5M5=?<e.FP3bU^@PX?6U;3X2DCY<:FRYVYGA/3K
4aaY;(\O250D_KCa]96UVFK8e^b:C2@.(:32OdJ.:0C,;c/Ic7gM/T]gUJ7(CP1T
FZ]L-1K(d?<+(4P:A#b6^^B>NSDbc+3/G-b:_533bWKWKKW:C05&88QC<[e#;LXC
^9J(Q[AUHS>P^fS+>HJQSXJAQ<UKK4]4/R1J2f32<.cOf]JSS;dQ>Jg/OPJP;^Sb
6(d-(V8ZT;(SY]=PCV:4\.2/ZVTgJ@e9858G&N#Q:@Q]]B]&gU>,;Q=MM[b29#Q3
LW3W\5O9#[TM>BKS<PG>#HB61fgZDfH<G#_80[5OYXXa)5<^>b0(PYTE;_&HDRF)
fIT8C45E@VgM1>c&6]C?88PK_:>Zb\aO?V,\e2FK)BN.#O))F@\F2DIT9_GZIE:F
.HF@:2[5FG4dc)8\H_2BJUTab<KDK,OT8S9G.:KT\0JL9c4)FHG+:D:(]>W4#.HN
E-RRB-f3:5cPFa,+/I;[&\D8-B_7JLM,<VJDHSV\g.1:.D81B\G2J/6B)UEGE4@2
Z>).X9+ffeY)fgc7.GWV#OH,4.4.I\U+7?RF6QTP<g00)4AN8WAKP75G[W^W?QbG
3I[7a,EOPE]]eK8>7ICNa#QP24C4@)AAM-)8ge973:\89cb[Y1^d(NWNBPe^@R5,
6,/;.;RO26&>Oa@6g^HMI5F6@4Y=;8VbPWPf?>GdUCTC;e(O;F+d&F.K10E<O6Ng
)/B8<>U.M4dOf+FY^K/c[,DW+E[g.A@J3265V>.U\1F.&ZRG2&R^O;JSGWgA#OH9
=-5e?K8?&_Bc3UHVD_d/HWd,Y7T:/Y:MfKC0O?@=K@.g_ARZXJ5d)>S6]A\=H5=7
)@PR2M)-eB/Y)YCQU4;[0=(Q(R8/P#0PY:QE&PD#6T_dWf3B)HA/D6eb9+JVTD;c
K+AdXS=&Q0A)38@38LUXRI<NLG1A8^N3.c-52aN9.+Ugd1AX:(:.C)TP[\)=S&6c
2:H&A]B)>1/4d>LC=P.1bIM;WZaSeM1cLA1D4&^-SL,POJLV\^LE3;PVY<@6g_<#
9DIFAV56?XJ#c<53QBCI</?SPL,&_(/gI=FYg/5,E<e.ZERD_Ha&SPQ>-8.gJ0]g
6Uae<cc3ZA9P0SAG3H,C7gg/.3@f:^a6AY1C?[MD_L5[_-7eV9bS&R)6BQPZdR,N
Z_V&3IKS^U)0H7]^5YOPE^ZLM-&-JO2\2f7&@,56Ld89-<U_G-J_:gO>&D;#X=W,
?JO]fE.-B;9@A/T1a,TR;8[U;ZPc>Z:\,&I-C]fb?<dG]#b2FR/=2YSTd/JZ^RU=
[V/BSK)SE4/[c-R=EB9/6N7CM)Za24HbLH42KXOOU>Og+(Z315a\?FF:6Ba9Y=Zf
EB40U,19Kd8[.A#+UaA^HfTQX-8#1H&PJS[ROXT=FU2QK.2eO^]U+e:U/S-B#Z[S
.,.ARCW_7?\?#/_=HI.HQ4OLWA_dYO:YaV?Z=XEIO+GMX2H.LNDTbc-a[OI1gAM2
fgMRW&Q9D#2/^MAV.Z:H?QB&H>F3,28FZPa28?1DL3Z/42(VL9M#5db]]gRL&eOT
&\b[I&1DE&MPS)-UN4F4CE]@,+59-[.>9KHEIJ?[_T8]W73P5baX?+><]6IE1865
8=)0><(2Z/ec>GX\\QZA;Od8bH7.:#X+Tb;ES@aV0DYf+61gA?Yb?>)b-S)dLSbL
(CUdZ361>Z&\;MQ+>Z3F09GW<JQ?e-]NEH(bXB,c5Z+(PE61K@=+YLB?FWUPR#AO
F6A.):9;Z/C4OMVSR6BG4_J#6N]]G&VPbTZ^1D.OPKDL>0a3H>[:+GWJA41GR_\N
d=f[K61L1Ye4O-8W^C3UeeIS1^IBCA+VT);Ag0-9U>bHf1Pac;b,+-gK;#\I<d:X
^Q5]DbXfeJSH>,/.8G>LP5=@Y)^a3&SYS?ODJ.B#D-6g975T):D=e,SA:.PFa1&+
F2PE9H.R5W.1E\e:E3PMH>(EV19CDWL]E13C^fE_C[:P6])B5W^EfZHSIcD<T.^Z
M@g#.(^@9THFS-.CGb93P7E.f1A0VJcfd2R1cN;Z=E602A&-)[)+PFP^b7bY?^^>
VU.(&@bB,@<[XZBF@B8\/?(<C5H-PaEYaP9Y7(JN7gI;1e6fH3cTS/9Z]P:_0<^:
3eNE7\VdgZDQ\BRLdNW,4D.:S&;?FW=S6E/3AF;(39;-^(VfgO8,cG2_LMDcU0#_
.@ZC+5W@1+DZ3G&0c)+P#GRcJNOQYSJAC#.PF:9?+3Y.=IZH\1U+^]OC-d2@?^-P
#:7IT)ZB#,)PR:<0[^751LKHOf@6AN@(a_a_1E=F[2TcE,gPbf6bWVG,W0/PQ<FH
7KYM+M1>JX7EG;0N/[=6Y4:D2^305cW2EE>N?E:.[Ya+40;J;5Hb_X9gSf&GT<T7
TOX(XY?dZT(c?2,[XH#.b5ZOf_H//f[<0ZI\(]DK07:H#X+Pg^Q/Z5Y#S;QW#&D.
Z.DW#35:NOV9)R7&@)fa9^K#QgOS&?(?0c2U0C8Eg0[J1XH+cN(\7U@c-aO=5845
4Lg52.Jb@g5G<#@N,U9VMdJO<>2H\5T-bS06eCZN3TMC77-L<<;2Ufa.B6Y)KJ+]
f94dV[/HA_?\AF_bGZ1SK8?(fdfE2#=PCe9gAXbS@TEW2V>-bU,V3gENCWAVUPb5
&fb_G2[K.+1Q<24+A)XC,CQE81H]\IF/N:J;61GLL=Ua;=2YXO<7dY^TZ:+)-(Cd
>H;HUZa(3=gZXJJ;b?G+EVd7A&V3.^/&:V(9/Y.gMdC&8fA&=ATMd&b)CZc:,+P_
/.Q0\^,(\1P,38K\&WZfH_f\?8XO7>M)ad;I@XS7]H=GAG1Z?48QO.#0<TJ9&4Q]
c#Q[0SY16>(a?=S2N)I@L.G0a\)Z/Jc&F7f#/g\:.D.;1P/D4P:NQf#8YX98(fe^
;bPXD5Cd9?C@,g1[7&KaF?GF(@bVQ.afd-8K(R^7]..3f;<dgf,MgNHGbf-&51@e
WcUR.8T,([5ZDZ)c/Ca2>^1HG)5D7W(:[d:fNMJWAN\HD+gJb1#g)0C[-BDg9(=K
4G9dAS[Hg[2(K_2fe/Ke=?PT@EP1OK6IJdGILY#NOY8/8[0.OY4?WWVb1657d0F9
.>MTOT&6>6<XT])4bJ1M@dCNXX&\<5V.2Iba2Y(UaC2O^><I5,H;8G/TEbH=-7JT
e/D2.^=a^965bP+d#R^)5,Pgb2AYATZ4B[\6Z_.EOZ,-[<FC)dbDUPB[IA^+AP)P
G=f(^>ZT)QI.0Y_OeF\9(EIb,:KOf2]\NcCH\D+H8&ZF+JZe]cW)II=(fK-^W,KW
.87)A0I(\]9Y)?d[NGZI>3(c0,-Ne<-7a9;OPOCQN(Q4:2[CB_G^+<ZLI-EHO\LZ
dAc^LQT\LY-Q18(MTePg;=aHK&(O0W-.6\_V=,?e(gfTTZY1/T,LfVa,V/\^aE=+
B4:+64;R9,0Vdf0KcG[a)cA8QR@2D8_L#\V?Kc:V)1BZCfDAB9J5fEGV4fG,G]KS
D08R4/f@BG#+57]L8MHd+?>5559PL+0Q\Z^RQZT5D]LW7-(G:<c)63@\]2V(;;YS
F2[cTb8O#)059?C07ccCJUPdQGb8a+3E(&Q6;=@&EQOP2f;3TcLL>CX@;&__g>=(
2X3/:b>XB)BRRP9D]K,5R[F[FGWF.)Q\><a3=[TYOfR=&VEI4\ca(aF+-OE:d.\g
I<#+A/),A2@?]W?>EK3CO>D^DM2ZKgJaQ;g(W5M+0@X+2=GHR(5&G_3]N6@8c)JU
.a54DO<(f5?6@X6H/9I9;3(fC0JgW,/H/[03g6T-WAT6gC5E[>ZH/A8#MYK=Q&&Z
c^SL<GCU8NQ^#UaH1UA..PCFV:M?KFLb90@-]813@GF#bWT[#gPH(S(<Ab9RH^N7
be-b&9JOO8\SdV#BLeR\F@BB)HACd[6dAJWf5PMIEP.H)HfD2,_c9g19TXSI=_#(
-:\Ec-+6I1DACMVe]gE:)ZMSHf28cBX#g[Y5)BHG_9Qd(\L_f(IF=1[@#>[dg7/E
(\g[M[E/?Q6IV@?L;;6G@MdC56A#D)-E+J-ID1VG.;bD_WFMQF29[L\<=XD7f-U(
&)\RBNX@516L.V9fLM1d8=8ab<B1Z4AZW-f+HaNOJJb3/32PYFIOTSBUdAU77JN&
,bZZRHb6_T91SQOE07BH,^03YT)@F50RG.5S,,/U#/fQ+Ta[<.?03<+Y(;Z5^6#Q
f.+Ce.88]J86SBLP5J:R\b0NY&<^/3..R=T\;b#IYLXFB.SF(e@7Q;0,J(8_P,E_
F-.+)<3]L/=ZWMCUU=IKR\((WgPA_\\_2QB@+dcOH:R5gUHdLT6\XQba^<JH??6(
=[&Q89Yd8,X6f:3a.[&FGba.4^1;=084RaAHY8&bHFVZ-O7QX^YK?ePE(K&C\#>8
FVOFKJYUR7-=+05<gW.2RELO8WP-1[N@X6D-<C^gOWOLeT1_RP[ML0:-1HB.R4Y0
^R4YP_2VYg.e;&5<UeHPBGVAFG8X7GH(Z,S3eI8V<A0NUMOJ<f1JQa.=5CYDY:>f
E#HW]H2)_JWT\#fcgdP6.,IG;a2G^U01Q,dJ=RG0)B27^GND<M@\T&>I@g6#6F&.
&AQ.J-VVUQ#G(ST+677X8M5ZfZ:He8a5)JI@(=[.d,;DdV)eVFE0/YdV)-3A)[T+
_]N0DW0Db2FVO]^9=Ig/VHBX=Kb^KJ8Y[fbdK/:eZ=)K7_O0O\T)C8W8d)1d^/8Y
KBBWb8E,T?fP0^EK3Id_46,C#TRUU=a394-e.TV&;LEYe^<E?3bN5HDK0^2adTM/
fPgI7Ra.&UXb7/=\B)T&@WSU)3:8ZQX#PV05->B,E7XaJ>X+-28C-3F&QdGZ?P9=
((C?/>.gUY<S&[14E@2)V/e(PHD+:^^:_GZUDI])1I2&dAXJ?0@EB4_^+L8U-XE=
AXbQLZMbJ;9Ne]W<I1@G&bGNXG9H>/O><;4L[:NG91SG.((]UNZ03;6RESQWZSTb
M/0O\:S28d+2S04N=\Md>5a7XM]fb7@L:.BNWL84._[Q2A@\;Z#IJ3EY5c3#IXJf
c4^D@&10K@I1A(;N-CL60:LeAW2@6?JY1\PBI__DBTC_ABY8KT#N[:?>G<dUXQZ-
bY:c)XCB._?GS;bf#ddXGN..^[=7QC@G&Y3FgQ[.FdC6bQOEbgNaL,6TKU]J6>-d
aAV2G0APC26S9Y9<C<1Y,QQ4/-<Ib4<MaZ3:BdNf+NVBFI[dFfTf(+dH@d<9cd</
UIK@A(UE8VB>CV?AS]#<F_C^L:]g?K&]R0-acb^W3)3IG),)8-OD4AfgY5_B05P(
2VbUJ)f6/JM,c\B.OO+)]=\,UbLOQNO+9SYf5;Ja;TP#d5H9K:[]6N40-AJXFg+.
Nb.P:W@VLXf3WaO?8GL5/);2Y5QA<HGT;M1eV#VSb:AE&dRcR)KLTFDW>#9IPCdD
Y,:4RUPPF)OL3\3YcA7ZO:CGG(=_ZGDM7a&Sa4VNT.]F\^1cT+EB6=_<d^,Gc=>f
d_RfP,HW^Y9E;<38Kb_2GBc=Hgf8.+e]UGH0.SO4(0P#BSU]bODd[74H_4IN[#Td
CMF9:ZW)^Y2>NJV?CJ_M&2.>V)4GNfJX(:W<68M<+cbK/+H&;GA[OWfRSZ@>Jag6
GSg-MU^D7@YKYS7H]a@fIR65@R#L7FA5RLM3c@^,)5N4^9\acaS1J[-L.dYW5_KQ
\Q>CQNMX1Ng/0QR8f)XSZ?YLbX.,;JdH]_5:KY>ZQC.C6A/53PERMcP.9IW2[f^C
S&5^FV>M5\G;VK#aN#VYVLU,S_55@OHKV6TS_Mg>>4S#5=#TK-c5]@Nd-QbFRcW4
fK;00/b.#FM92K<J:_@/OJgXC^=^0&D=^HMUYa6Qe:42DK/P0INTTQG\T\IBf;Ha
@K;MgTDa54aab,Ze#GA&D//[?C&?@N2f]CCFe;42=4+GgRM+K8]Q#I,V9C(,W0\1
U&L-??TURaJcQ/G6b<;R]+b=+@B:Ded5NY)/ZZ7Z+CSe&05OP7f?1;b]@67Ig0NW
GTg6cWL\66cIAf\4_W;ZIBZBSQPS8cfQ\NceTK+H8Y2<?E.gEJd-5SMLCCUOOUP/
(^HBKUDR8<?EaPC>I>_9)PZY4bVdPa4/\U(>_]V_,8/P2\DNa(#(HO9?9P\c;I:\
+e+JMQYTbg,/,YS7NUd)fZ[f-OfJJ8Gb>AZJ>]3.Pg10\H>#X7M\,,HbBdaHHg8S
/6&GEL^,3BVP8+aAVX498E=42KB[Y25XZ^DW;O\9bX@^>^g57(a02LO7g>e0b>IM
:0BQ^7g+?EfedC>aH87Of1]5[V3J<6JHGZDcJ:@Y@5<,PQFD>KN[(@^cW#9K=_.A
bY&O3<G\T.(<1/39>9+KU(bPW#[R_5]K@Hg/?1,6AB@?Jf^bE3d93<2]Ke>R2GMX
DRM3J6,B5MHH_JCV2a0K,-C<gU>SD:P.CC[gDZCST;.IaUHJ?[+0IKV5NNA(+H]0
DM+GV,I#Q>#N6I;NcFGd3T;@[-P<TR_16].gKVFV@E:Q]fZ0R_AdI]FbGQ_-[4:8
WdA4EgGMdRP-1JB=ZV-@XFP&6N\Y\<@Hb]BZ1J,T[OB\c-7:2a8+b#K#]CI]W0C5
L@CLNP+(,1?[)^V<TWX([KYXQ=U4c.M.]T)2=0#<+^BOSK8UfHD4I,e+RNWN\6WP
Z&Og#Ae;ef(XL2-5Ag3L:AG=;#M5@<[,11M:O]Ve(33>2fSP.(H#8@9&9N@2?R[5
GAN54XRZcU#C=1JYZ(8BTRTROb?F+>g)TTU)#fGJ/7Z;/1\_7?ASM^9bJ_Y8WK^d
a+5dBL.:UR,4(Y9JWF#.+&\PAQF@gG1F12fMGSdL,ffGM#V.eUGVXC^66]<D,3K(
EMS]7dO3)<?LIF5OJ(K5C+KT@d)<2(f;2#,-R4ac@YeOffF\[V=J[D.QHSgee4d8
P?V_X4Sfb10eH;[VA[c0RgP@,@@XF_RYWDT=.2Cd0A]bSMW5UDH,\^M;E.ET?S=_
cfA^+8W[H#0]A;G]UTf]3H(2dSN[GAg_[UJQJY83[BF#fUU/>BU_-D<aUG2A4<Y7
U>]-9RNd),ST]g1J?TDB)GH8BE8&.d[TCV4_9:ZIQ7W8&\#FGNMAbXd;:^_4)]H&
3]D\7#?,BVIF<:\/>^\(WWAAMRMP0c86BIUd?c)aA)3XEdO::O#ad8TEV-K2eXN#
CQ3MM8QE-7K41CXM,.WA]>P_5&<_UI=G3/YR5_(#0LgI(_,BGG[YeBa7<N-d#e+-
V\7^1Q?LRgH+_8Cd;1f?/cbK+5EeV/<M0T>,a4F?9CM&6BW5XC5feN9#8__N5F/V
A7)0G@W];ECIc.IdZBOA_g92G.2)ZR[WR5(,36Vge0GLP:>O8<6/WFJK56_YNYY9
eFRT=>Ad\T^QZ=?ae#Kf@;<;F7Y9?+55/SR6Ca?;NGVLLZOF+-?&E=PV8SGd_SBK
2FfXb][ON5LS23eSW@)OBEY^8A,#7ZFYFK-4#gZZ8-L5;:(NE9HbA8YA6XCIQaZ4
^Q?^:@Oe4A,V9/^JB_+@<\c.WMIX<&C#0[VECKQMN^0HD;K:X01:Da2XL^-fa[JP
]MO27)@=2F1IWW(+M<L?g;\7.E(/cJHg\=Z(#UOD;/W-0/>A3gd>?(\NV..5b<75
J>&1X5.JIbaM8EO^aY@[cWXU_NBfb9JI&I.W&1;FYU@3[e1C;<C7cMAbWdFH_<4P
GI&Q40BLWT5<dUI>1gKCD7B7]&C[_SOM&[:a)f[P##Ia_#RH1f1<8KXfQY[+(S;)
]SBL9R-RN\(4<)M@OOgEf9SgWcFQD^7UH<;@<72UUWHM^78\,,H,Bcb3bS@bA-UP
Q?8)4)MPXVC^LL(=:25FZRX>]BaQ.?^#IKCY9M^ETf5Z+4Q]e;NBLd)QM8PU@>FJ
gQOc/;TN[Wb.^70/5Oa[R,7QDbg<+)6^MZ0bZB_H,S.,7BR/\&XV+DWLB=ac)\3Z
L\dBZcaVCa[P6JAdX976DGN,KU9.3YE[?:GeF4OGL4],0VXW0[gQfDc@g8N/3[EU
#1YCQb&5MAL^Q[c8VE#S.f\N5(1;N5U7PL-]^ES]aB42^J+G8V?GdC#[+;7GE1?.
fTUA/RM-\bKdPVg^-H]9bfE>G&IcQM9&^b:#fN0-URH4H)6)PNcN-;NP&VDDFe<I
BHd<W6AVE<[C^f@aaC;(gg&cP/H6##M-U^E-TA2Cc@91;GRZc=ME@d7Yc6?]PFdB
G4;-U>aM=<FeDASLU/AW^U&ZI\Y[S15gEQ>NC:Lc\)P[=/]D)Z)P?a<c;f#^=2NO
9=/86<KTHSP^,fM_N/WWedeEc.cJSD?TF=Ra9]8WJ.E#17=7R38FHZ@GGMe@?X&J
a+(H1P(W5ZIaQ:b,M:TM4MW5c@9JaPVYd>#6,;\K1IaKUC5N]0P>BN@DYORSDO95
Y.PB]HP_X3gcC.:Xa<<;]_S&?/O)-aGB\XgbcB\JH2-7PE,<LRG5<UcMVVBOXS+N
V2UFYN=/J6b_9HVCBf5+W_aLO]:#F<b?C0^UEN_Q&1VWD/@RRKVFScE?^Md=\cN(
IUZV#+/:)ROFV=BS@@2@e4Z+O:NdH/:<T9R:Ea?80N2V6&(.K<^b]d#GIae];A:1
1<@_b?d?;(TZ#C(ZC(1^#)E(:>_NN@.D:@G(51aCcI;_LT6NF]BZX.8:KWb<\NVR
7TeF)=/DM@e45Q8dR(c/c/X;A]C12?8XC_EedJY7fMUM@LM=NP3@G66Z7O:0..UY
NLg0g?.a>^6UMVa;.GdS^+b-]Vf\CDfTUENe=YfYGJDE)@W;UJE]>\BF>DRaF3V;
c7CELR03G_6M:4XWGf-RX#b-aeSZ[OYWg)QA8aYL>M+2eE)\5b1g,DF3b,D.S+.>
>9>CY./DV.FB2(d2K?,<cT#N=ZIdTHDR>(]fBYT45ZN61KZO61JDObH:M96bG8GO
QVe?,]^UO+O\gY^3dUfA)>HR[ZW>UYVBY-A;3a\L7+=LKb+O1fV4d1c=>17P0^=Q
SGa@HDX<&B=O,c#(4#Ia37>2LK;&L_c5D#]5aFed[[+&M=9JP+BS&/e51E3IVV<B
;W&(Z5BV4M<C=WQ01M/5M]15Te,-ac4YTL0cS)SM4eM(06RF^<JV)C-UR>DZIY-)
S&=4.Fg8&82&1U@])<VdEVBdJ96E-OO[F#+/Y1SH[HNY+>6^#<:D6cUT03+W8]A7
C0]CJ\4-cbF3g#c7;,@H?UGB?R<BJb+K8(>37:DC-+PI)U_\O1U+]f[C-bPX5K.3
;O(X\<c>-3JV;C^M-J<NAY&B4.6@1-LPf+]KDg^K;PTEOYR_N25PR4_0d<Y+@cc^
N3S]((DS6fc?T5):(7@^OJ@N#,V@G7\)gUaWfR_)+A[0YBdMCI0WR46R?EeA_I]Q
f8X4Y^bV)@(/-/=DN0b^,#;^48F)_ePT,(G=F:U.CGZ?aVZ&/,#/Y/HKC[E<5?cQ
HdQ&/#FFH54&1[1a7?eT2e.Q-JD2^<MaDdM&^F)>+C)a,g557JLXVP/#F-J1BPB3
\))g&)Qd&AV2GOP,L./84M02=+fK=E.ST_)IbJ7@>2cb&SF1JNLX+YDD>TeIgC/-
,1U<;GC2:+(a())0-WWaS@63@@N_=QSR[T+?Eg2>]4bbaJb0YWRZ<LUI9S)NAc[(
^MLZ1,V?5-:6@JOa(e[S9K\C[UVJIg[)@dT>,P#+=@L)NV:eP=WYC8>/1N7Pea2E
]#KV4F7d/Pa/K5R(&.6J4SQ8]JG-RPEU^Ub.c\J^+<Q:J5b3)QQ,Ha1If0LbI;>D
O@+&,#O;8LSH=?1Ja[S,5<_NQHB537RUALAJ;<;L2Q;:GYY3VEf<Bc8R\YO1?dGU
1P9P)DZZaTMdHGXBD_V6=f1?3QgIIDPS=X6-(TZ[f8N]O6bV72^<bR0J5VHKf1#1
^3GUaNe7e4d3Of\>G_KIT#UEX[/9T)b+M-/ZJ26efHAd23,^,VN6T9)G3eS:OGNc
P#[8Y&GX3Rg:TfN1-Q0<&PXV)L&.d\=:W@EYY7XQ.D)948T<HGGN@=G=e659T(?&
eD0ARTO&c5Xb4PTXJdc7g=F_XaNJ84>&^Bd=HOgJ-BcYK8489XHc8.^<39e.K6>6
Z[_X0_a\3);/]>/f3(XfAP6O]IWNgUdSZd4a8/3=.^GbHd^;dX5UMMQMJddc3+XW
.<e(77^_/D8aCO#::+T9#KM]6I_YGHg,L3NZQaD]0\QF.gMKJ=.YdJ7d<4g<-0R-
=LbGY7N5;P873Da]Y+61UVY6;-OYJFK1W0B)VRfHQ?0c@0IFQ/L.+WKG[N9ZH1-b
76dFEN_Y2CW7LAdTU/L)Jg>4\SX.cP[6@&I^H09G:2&ecd/=7U^g8):(d94DA=Qe
,\_3ad6+;\6@.E;C^1R&d(M&+\OI070ZT8bQI9bLX_EH2Q5-/f;RC=)=QEP4X,7K
J5<&MaI#DZJ)@XTZW:WK[:VPLdW,=C[J&S>TO)WbEOZ&>3\_633L6R\PD>Y.,854
-U]e/CS7;QZHdKaEC#>>0V.f@Vf].Q@Z&C__<_Z4>N[<f1e>FO>JEURecgCP#9YG
\O#<Gb-TcGCMMEA<N3AR74^Y?2-Oe,&5U;+JV=@Qe77R&fUXT2KT[0Y9]9.-Y3TQ
T,Oe)TGeTSbGdHQBUI4H_QWNR;..R&(-&3C-5/PQB/Q2[UJSRS/?-dc;dM?^E-1=
ORIXY?D9]KE?@ODM,\aL0^4U/HW,UBRFO4N::@OD..a;bf04B(+dG05,D-6,@Ia,
UNFb6S/E;d]geg=e5YabV\0D,bUPB:,WQKAS#SPZ:HVI>Na48_Ee#VM64@c]A=PJ
T1>b.T75RWbN7G^4?&BU/P3.cNO;aZ=7[aF^+8UIT;5]TfV-Q1>N&/Te.,[=^A2\
8ZDR^(A]H&L,e#KHfWZ:X^24.TJ,Fee=[c.Y7&3bMS,SK)E+.Aea10ZF,(+ZMN^J
:HcNQ/V)HbFMV#5EcJfS49gS2X=P]2#@]KDb35O@\>+7U>@V24CceS#ggc,\?d[A
H;g:.a7BM@33d+)^YEIIY5O>a82O#SGTG7c_fXL?N.Ig\0#Z9^[.RDKQWTeKdY.;
^>#K2-6WH_H9-e3_Sa6?SFJD?b[Ka0d5ZRJA),Z\I8c4,3(;K)K=d(TeW(SLBFVU
8)^JB\DBb)W6?)X]RA>@?MD;2PO5G(ZK<cK7Z47>NIXR&PfHZ;EBXZDY_AJB)G0H
(BY,XfX_+IVL9)PbS(7:8WBY4)DL;K+W6>\RCK045;d)C(K25cJ1L3-MG\GTH>-c
GJaJ+)gT6JXW)<L?UZZ:B//NW/2&85Yg[;HJU5_#+JDGX_&dLQ-)?@3ZW3C4KQN2
c7edg.63]_Y<N[\<UMQcV@T:E^2C<-P[N^@_SYBZE]P:-9S.g_>gQ@#\<Pe21IXN
_SAV02IR/ZL0O2VV5N7/dV&1gYRdRH:H@]PWLBA;M,?O_)a4eDeT6L6fH6_&A+K^
NGUM_^B@cc8@XUU8)PGZSc>ZU9]R;fe8TZ1(8RQCb+:]5_/XLd4beDS_EL).SX]H
UBHHZ]^&e+>T&We0:L:)9P:,[ZV3URbfV&+aTHUINgJM,8VA)955IAT[92=-SM5<
))(Oe:3cOCT_N@_FZ8f[YA.^XVG:PP_E#0HZ^-g@0d98NXa<_g2F,bYVS@#2cVU-
^WEDM.7SB0[UB;KTF]MM.(=N5/fGLBEd3?IO#,7PMRXO?C2KQQ+2S5\LC@\MA-N1
)dN)[0E?4MJd6b0/G,V[U4#Mg9O&EWG+b7FgI,@NB<DaG5\A?RK0gS8+PIf(P2WP
VORZA:[5]7Ac>SN^b&63^4\<2KcP.f.DC#Qbd]NfP/P9PB2:+O/6Rb9b8Vb(fB>J
</W@N9/1KR)f8VN7PN4U(GJCH+#TS2\/<-<W_+^[(XR\+_\(LVD?Yg\-Xb5G-<(Y
)bG)S>/E?W#ea10M9=B)UUI[8WEJ.&#2\Q_-#\]=fQ()Yf[5BbH^#5.M3K\(C]^U
d./9Fb.M+-P]\)\H[PI[@?g;:J3-A5ZOD;1<Q:2Y&S;YFHAa;D5B=@9bbLC)]:#)
?Z)gQ#9RF,CJ>.e@X-ADIDG6ee>MK.)?UQL+a[SVRPb#?],XS+CX5E:-ZQZOJK=M
?@cKEU5N3FM#X&R,>,EDaN\@BV;f0g3aYQgPbIQ-;b&X84,1C]P5P17Va@bA<=3N
9/8g<QX&/Ef6TfXCGA\&.,:L-Y<9--=@Y(V^WMHCZcSS0R:#_YGTFMP&MdXU>L&:
/CB]^_\deY]&2=Zf:]0-<.D)Q]H(T0A6WX<3?,<41?eHIA>-<NCJ8^67ZJ[?S&8^
;@g1YY2R-QB?VD#_ZV;&H/>,C_YKW9cO]6T@bYf,B8QMT6F82/4C#;^8Zc-N5P3)
-5G;TV9;M+>F8/VJdNDd]GfS+ea0^;SOb9W<LHMK-F<)V=I]9:53L9>:LZ1VH>E,
NI&9fJ(I3gIY#)8/]0(6_&U0+D_[9.D:4;M7b2Rc<WCJeFdfG^V1I9_^2YM&6&0-
JUd&IbTNP\(4LbUWGKJ?_,XTU8TV1)\-/5G<],Ye-bMc;V^:(/:cd_(46M6[PX=>
](1P^2_83/]FPLI#d9ZWW64(JMd+E9ZM-JUS6:P^/a&O3FWS5Wa.4<@G.W^Y<+B)
M+(:;\0TNdUCQ]ST.,N8[6f5(M]Pca969V5T@<017A.YBEJ4c]FN@f.8H616aEHc
2T]G\)L^EU(=6I1Z0YV#6:<d-e_@(W&^41;L(.5:,7]M?-<cFgb92g&?>J.f0VME
K;0XI^6JCZJ9g7WF:E6._;dH)F1Y+dPZ4db>O;Jd&8KBY>FTZd:BQ[.UP7(#=^YB
UB?(^/W9bJH@/&UIHc_[4UJ<b]>@-3T=OYce3E52/,bfN+dg(\XR]@\,d?db7GR2
Y+>d(9f-JR@AUb6dZGb,cCg->Z2CEV/M5g?)05#F6.e/)NMEg<E&(Q(-e]>J5bH/
RZCB)@M_HX>e2SI/.dOdH]&+V#@731D<b)OY&>aAB;8:M8f_\K22QL-2f#UbDXMI
1JDY9B(V[KeO3=M06,63--+bFSVJXF=D62WRO(0W)G_LaN-\\ca9&I1OD28Z;0>4
.&3_I=H0_4ecH:N0@NI#gVM;3fcJ8N/B#4aLID20X^^7UN<g>FgD,ULR:64D9eaN
E_4Y>89BTJY:;B4\f<@^P=OAa;N[OP=gH1W1WLQ;HV]GB=JA=#PJ\baTFS_GbQ[B
P]>,HaC[cRB8^XQK^WC>XOY\.b]J,@8fK85a+.+Hg\c]D7SRFWIUAd,EOdYf#).9
9WK9SN,X-U7W/bJ6QeddB)S,#XHN/:=)WGA[<J./+6P03TTYdO]5>@Gd/>[b3^\^
a;ZSY.aD\Q[BRDG7eeK&CQbQ\Wb,1)XT)4YF0Mf/Qf5VM+O?PA](\?bMLI6MMP=8
)4B<8:FMXI9>ILLL(dCM,d)>^G[g_Z(^g.-CBOJY&<P:EC?N6+J3f<]QQ]@c9LgU
8YT=g0OSK,H(R#[+c2ZO96[ebe350,XGfER\eBH5^cLY+DDcP0IGC/Ng^\1Lc=X\
Lg<)?g[4]DV2FQ1^LA^SS40AK6Y2D+X;JS.&-^0fLRBYbTf\[BJ&\^dS_8-TgfFd
G#]O)]ADW\6^MQP-@2./5S)4LB_[B?VC-Vb+<4g(Rd5O->SFHNO..NX1I<&#F8I(
)^)).+[f3=MZ,J6GPb+d/b)+F2=IM[eYd?49UKNc_++-HL/^;9IEKdb=SVdF_<KI
(dAP0MG_<a&E?M]=:78L/@6@NS9D;NE\c3,OCO?R>CXB_-Y4[4<#Jg2+e6]dY\JM
B-S]V?+c;7D1>VfLX0-=:47H8?WDQaVHa,JL]:/PYSBR?=;<6B<0B6)F5(g^Ge8[
6JP9bV]J^PT:5PD(V\g\VBV+KO/0,=.<Y38X-IOF)RKQ<<W_9NW(6IZa7(>M_ICD
;?76JabV(3JEWT2cGG5e4R5FX/E6OZ\,0EHTg&[5^5D.=LZc70f\eTa[G;9efaQ7
(5;.V],cD=[-g[9XZAR7fS>ZeY#aV1^[XfZ?)F3K<V@F=AB#e:KZ2bQZG^J#\4dW
5A-<H+P6Ucf8Za/1#ZVW231PcLCV1L7c2&@>LY33g<\b54,M6I3&<CL8U6d;B2cV
YHOgGZ\;YD/,\Z3_&,f-T37QgX#QPFFe61OVZ-=Y;G^5I5HXIWd:NC\c.9I_)E1=
OT6cX;,RG#b\c5gU\?2,K6G#I4IECZ[P/g#]RbWMe(QHT[F-bcHWNa]SLHSUR[]0
0b\XMI.cKJ^&M,#)gMG>>9FU]M[ZJIe7BEfZ^XT&Sb6_MW?W.7?P\DJIPBJFA=6&
R(J&]aE>CCO9D,6Bgc_\PeH^Vg0)B[),9&3Y(C4F\M.&#\fTM8/cP71b;)7;D0I(
F;<c@C?OU1ObXO>P4FG0a\b[8]&gG><6b(/aU//QC;OdW2[WLBea2)QC(K6Da9Vc
\H.WFdY^\6BR>.B;?P.N1^?02FYZVS,9cJVB.^XegB^Oa9AUX.W9I\D\SJ1D-4.,
c/WBcFc#S&Ld.9@^gDDgb6MU0;ZXV8@OQ--K<^V22&98RK;<X5cfdTKR_Vd>+6VJ
<UL4WFK2N9XG(M)e&=[6.W>2W:3S<733_FHc<=@,)LW81^\RGC1W2U4@XOT90f?Q
O:c=dUXV?S,P]gC]NPfZbB(\8(&gZZ1d>?P=fMXXWOa)_6(L2/cFQS)[\aUOeOdT
FN)-@WQ7.CaL7CMGZJGKZ3FA#:JN./B<aL6O54R0A[7Ng_C\dI.2X1[7@,T--9WG
4X6?D[B@c)H-,M+ecX77OSW<gX4&VOTV>26gN07[&SIbbLfNgBF/X[M>^O>RaY5,
ca3;)<X4N6T03OUU)G?=7]OPDZNS94EWR^Q;K28UA-77>,8QV^X1]&Ag\?Ua[FGd
AX1;Y2GdUP&@N[YF,f\48-,J2eF]T6GR)5]\_72+eI5_F.V)eO-SY556VXEAL/.Y
U1.9>6+I<fIIgSb-U7ffCTNTY[]\[=[Wd.^S+OJ7M@HD[f>dIM?@8f^M:XM(99Ob
X_P[9#dF7BHHN^:YV-_(5Ya4AbC>If60Q[U;\P(LA[)]XJZG7N+##.-<f><ZNPOT
^,?/>8Uf5aQX1?WD>?QfKTAHU&WN(K:LBDW4?Q?>@#TPCUOD2AQC?T&:#TR<R92]
)G8@^QS3D.U\QWJY80Kf6RcT(B=&3[Pa8VGYPSLNML<KE]CXTCPg5L.\,8Q9JcHW
&JBe7BY5]BTb4+K+)=4Y^ARXDSOc25>R+e=BIWJF<<57Y[dgNN18LF#g(RTG/M?6
/4JXQ[CVI60ELH:f[f29C4K9A025)8YX0FFK7=:;Yg?(/,+E2G23C6P4Q)O7eR[.
5ENJ.)1d5=ZD^);\4NN1^GQ--_d;F&:dC]_4dR:/Eg2KP2(<MWe_\ded</fZ<b:6
b:L-ON(V^VbZYQ]eE,QAQfPC[YL,Z4NND+Sa2E@P>(D?GTB@Z.E_Dc4aIV+KPaJD
>2X)AAc]^NGQBMU>Q>]9dGgQ(>OU+NN/e94ZAEc681b?);DF\cgWT^>\D]7+9+>L
JK#dESY_LQAQ4A<_C=U9e<245FdgO]&>==Q22AL8;3gDAAGTG7<P;2I>6MeS[RO,
/?IKE8HX\GZX8fT6EBW3:Fge2UZK7<UXf]LS.-83];EATWgIP=NNcB<<NZ^3f,RD
T-+a.P6F(d=NC3SG;P+U2P/4HfYP=X)GNM:@MGE_6@M7:V_Y/0B6/07;9&_IU#9H
AIf3CT]V3a=_8+U2)#LNF/fELYdX[Ea.(9e4LMQ8I+F^4XD,5IAFTK19U?CJD4a7
RWT<D_>QL&A&]#(>XA:7HHK:^8ZD-CBXZS\;FYUT^0[8BAcDFW)MF\/K2]-_;_aU
ggD/.EUW#AR7+SUWH^UKEN>=U@Dd(4,H:7TZZG:HH_GfV[^?[HMg<;7H>JT,H9(D
OBRT>Q+[;BIJPFQW2g5E;gPZ6))F?<I[7fP_ECEIK_A>-6:+32S?5?4NJBTRYZ:C
[Y9G?E7L7;3B,@VOEWU5J3\#RKMAO?>afNCa_8S5TO48YU6C79.J#D@1WDfL999D
R?49K57,7>&09IJ?c@+eM=\bL2+,f_]E<\?L3)=16fZW@57.\[Rf&D6e).c>Z,;7
:24M[GWcAGdE)I1(c8dgFdb?ddE9f4OTEXLO52Bc4eP,H<[3E;\8]O[F\L1>2@)6
S^Ze1WHbX?3>ZHV42TSYKI\(gfTfWP(0Q3bQgZW9.(Q5A&5F[>V=]27_T6[ZeC.T
X\e1D<)]_Zb.=#^@;15NNKDde9(OO2)SL?UDVRb:/WbK=\O.(d5aY2N+/Q8<O=98
PI/]Q<:@[.I29?=a,aR?:>0I/X^0@@g@27F?EN:V<e?g=8:C+=NU=G(&90)FBG\A
\^<c#3Q9LIERe(S=Va5?Hf0:b30S_CfMCUbe9+#[&01cdYM)VA1JB[gCI.MSL4)2
PVO5KO:B?C2791R_FcJPDCb-2N&QYZ^BXOf&&RT>YGLAYRb?4OMRA&S(271WY()A
M\A=bW0eOB&THeg7>A3a39aaE^[HIF(]FLA)W.3[ea.6YNF\C7_TL@_=&5R,Pba;
]D&a909bYfF+;O+97XZL&,@d\VPL9a]P&3Yg9/K&T/ABIX=]ET.O=C:[?Y#.T_R5
M:3;E@<&660R3:](HBD@KCC^:)3TLCfF;E4[^(JP-FbWec[\WNN+E?1E)d]aW7(Z
=\DN=[,^:RbS?Z1dUd2VMUCD0VZ-FO#^9WGPg17?<]C1\8PgQBf4Qbe^:7BZ,5JA
PcFg9@G3d0)WS^;<6V5B:f1&7N6Yd\,Y)#M9-^DI\GP9@46R&bEK)9\)eN\J?XS\
d1B#=aRUB\[C-)TQV3&c\4>R>a#/eTGAI:V)JTC93W+ACZ)+P1bT/-@UJ.FM^P]9
I_7d4JGFP.7[,XRR/HBGEc+EB6eVCc[8<[UH)KDd6S)0DgYZV,L2)U1bLDPN=ST#
[DS7U]R<E,Pa_03a?G3bbC/6,aU:B=S<K:EeB;7=?M72a>Ze0J/c9(XeUX.gB]H3
8;.bRSBfT1XB?H^V;R<[Y80_bR8GcY/V9A+YG+^9?=E-a:B>YI73YV(==R.8HW.<
9#R51ePBI=LIRS,L90FT2e?0\cR@=^S1:?[6a#V@)I=FO0B_\bU=[TAA+[OJ;NV9
J=gdP1#\NP/D3#ZLYRG9X8SY.BKPU\Gd;-JP^W-]^U287b5.aT_gQaW]OF.TBI^:
@?6fMIFXSZ[(V8;VY12OEXIQF3BKDGI]_JMR,G@eX1Mc8K_^WM271.(E#AS^WCeC
W0(?9Oe:D1RT+3XQ#^(X5BX0]5CKC-\^Ed=bRON<KQNPBKV#g(EOT>5S&#C6?N.&
9U\aU:K9EC,f1RHJ6HO=2Q(N9VUATb3CQW81gdNadV=](U)U7K99ZV?Z9DUL5D3a
G5\@b)J)&1V,9c8bCV0gGA7<@#.ZT_I9Z:UaY_V\MCbdZMCKPGb3_J[fP47/dg,7
46f3JZAN-2H)F,WUTA&5A7YMM,S:&eV[[-FHGRd/Y9=dJ+/g7(I)_\WTL;g=1[U\
)WfR\-8V=:b=[SMAQ7CZ9#c#,+Z+7W5W(,UB(6&:JVN?MC(D1/CO3]XFV>&R2/0@
=a[ea9O?-Y,XK4QN.&PIQW40O[\aZP+<K:>/TM.(36I_=@,R#_T2BT2=+8I=YO=A
W0Z:?1^,ddb82CPQ/+ARI2^De+[fP57AP-MFQ61T>>-_A#aJ-F4:V6UeN5VRJY3)
YFZ,6R?egPILGa+I3:JT&)/3.Ra,:@J7F2Z@_BAUPD6&F5@gU..>YT+GY=?J?;^8
#BT,H@>\)4a=0>ZYe^+#R0TA9WX4;ZI7@315b\R+<.GRS4Ne_Y[7]V(LH@D5D9A(
+.4LTTa3ccIRXa#=0dXG-KCUYd6-3A5,A.DY,JHF<;g.HKC/aXN>QYSba_NgHW;W
;Y:>L(D^1[\6/N?dZH)OE2S^I)H@)4_H8_0V094g4b@:0+XI;/_^V)8INUQ4[3^H
&Wd6T^G</B83EQLG__O]?W6H7JF+@+Me,,OWdK&Ef8I=B]<c>RTR(e0X.29?+M9?
FDE-_4[(+46O2QC@d><9FgVQ&d\VZfHf9Z.5.7/B-f/J?.WI^J>;HGMA/8LU@Yd;
^Gc5A-?GYD4e&(_U=+(IR@[L#ad6d/S@9G#a./>QJ;4,A/2XY0R@EgfPA<E@4]9K
IA(c_B_M@:Z&)1AU3>_=+UJ9]De/.4:g_][g3L=/,S?(>4@5MYRDWgId+aNI[T0g
])=TG=[MFObM&7N:<TbPTLW)X=9DT]Z5<GaIaQ0+;+4bca]b^Z],K4HWJM:@N=S2
B73cTDYK@Z?]LJGT_E<(C0#e>\\<\_SKK14D3X7DKd#L,g^2V)5J-0A#7&D0?eL3
L#<#CV8WKg^H50989A9Ne-^f;C,R2RR>[XR_c>W5.L\#&34Qe6N(^O/K=g8W_U9@
,FSUSVW9::ZfdV&SE79F4MJQY2:(C^+4H&EX2JbOG()c_;Z5+/SKUZ29CET88RU<
ES\K-FU:H8_d4e>JA76#[@/16R^Tb-[-CJF2eKD.XP>I2#LDNK/.3=39ZL82c3-R
I<D3,RE#fPAXQ@N?+5S09/1Ga;,Y4+B,&J=JafXac)Qb;NM_H:,FC=\4JcK;ULRe
c(KK:3e3gP@&QfP:,J4K./a5Ub5SE==X&@9>HVd/Mg&W@HBD=0IRN<KK0G?EB>&9
CQeRK1;GFI:(CR4CFFceKQ5_Q3J]B##ZN#adY13-.bc&S4a^^2[^=_ZZR<8??0,_
DS.0J]]);L2?&bP)+?;\UTDde1J1PH2aG,PU@=UZdDO\=PL(5SYYHbO73e32Z8D:
g;MMCF.#;&&YC##,^2CQ0I-LQ]1Z)O>V:Yd8bXV?RSGY1I)NT7XCK>=/OK^89XP>
7dg0cfX[H;SQ(K3b35S623AEV^f0FCHDJ/1A@2&2a^]cM_N\K5Ieb/JcK;gX_SBK
fLRH5J_g9Wc>.b)H)3e6CTbNOFXU=;]:01eA\a2@e<K>7&BJ/+-Rg-EdPS6Z^ac8
gU#V=\F@OMgQK.A[=a>]+aU00-_Zac5-,N#FS6296_[E]57BU5?1N:.FO&ZFSG)K
3Wd662>\Y#F&fdK\^R<].0]d:@;R7WSM\ef=1;#Q[gY4:,,ZcbD.>8.&D,1Q0X]\
;A^;DP\D@UQD#VbG-U6IO\+GGI++U#\<ZGJ1+ESL47PJ9GT#66;GbEfT77ZN^MF]
JJ<MMP7NQY^2-20K+]4M5P\6Ab2S;F:8\RUO735Ug=cd,I_@R0=@Udb-<1XS59>]
24#3X&]7MNZ+b.TNBb3#(Za&VL&]V1WQ=-(Y;D=&07e.@BI81dRR0L8a2a6[.&+T
5RBFGAe^4::9-g#;2:b;VUWGKDP_K,?AO-^HS-MN=f0KKR9_E0Ab1]\-DZ=-4;0Z
7UNT?LcZDDW4U_D0L)/d?:-=g<4SLY<B2KWE+1T833<>?J(EQTT#7b-QY5;75SJM
\ZdY.f=MB21MTV6M#WW?YcSdNH3eU0c2CY27UZC:7&^[3K,N]H<AX/]T4KO2=5W1
V\^D0>:.G\M?dT_#SK5^&Cc9KDA-/H>Q-4L_WO7M))Hc22?48YgKPMe4K\6b_O,P
c\XL_M4+27/G5;1#_dHBV>H;a30b4NSJC?f-7Z8ga)36X\^.g6ES^)#P=YA/Pg1>
4b-I5],^IC.3?P64PI:;YM)Ne>FIYZNNP&FAMI@6>dQ<XJO/cY^[[,B2?<7aAVRe
AO)PY=#BT1(Y)VgeX3DY7cCL;+6e4PI;#WOBR4<J=CKB>.=-GC76<^IEZG?9G3>1
NM+\7b?3#eBY\0_e)J6_1.AJ.>IW;]G&]?b)2fER:U#eH2J/#911,>9e2<;5N[Fg
_bgOE6U7Q5U[0<,QDO?W7EJ=M97;]&Z>>UW@g/Ac7@/2,e8KfPR4Zd^@+(-I-\O6
@1N\eO5;QNeG=,c#aRR38WfAKYSe0@GX.SFN34;Ab2.)E2UXZ:OILWVU?/8C+BYM
g1>2F/8_aKc-B-?g5fJ&168(8+DY:#DJ@1/]g[(NT=PGSDPRQ/?\49N.)G=gL.NN
\Y_+[CN;DH)Y8&\J/B4DcYMGD=Z_e\+aV2IYNSU-]])b5ZA]d(dFV1Gf/bS4:Ef:
:VeB,)P1ca0,BT0;8N&\\1UA9+K<I,N9EZBAB:=T4K>LQSJ/AEMeG=+)@V?.2b34
Gdg^K,K<;5A2/A&@2T13PcdU,AJ3ZKW#a1E>30>:8WcW;LT8=(]>4A3FL:)dJ;XL
KYG14+,M.]?_,V8^GTZ@N5G7/d[f5YVS)-(^]O6aGd2IZJ.DR\1<JWC68gE(\)<T
g^OH\.Rbe#1.49RF2?LY0PfH@DV:9dHYE@):aR)BH^6/NUe/\8LSV.?2E?I??HDT
cALdICBd+4)3d]13.?&U[W1IWO[X@74aL;P=KUQb<.BK7\@)fW:35QJ)QA,B)\,Q
_7[<V]@VUFANLT_EY]FGH#[#WL#ZIE;^BQ9/_BVT>9?@D9=XHZGNZ&_@#cT.DB?,
>WAF]VdAJ=#<)4&>1G.>O0ZGOZ=OU-]AbAH<-EP=+T\VSDI<X/[>W^;24C\3_HWB
c?3eC#B\f,NL1gUXBGab7/aNC)-=JF1BVU07@^]SHd2YeWOCd6]bH8A7=F]NL8TM
-S:FgcV)M9f[X^(+_)Ce(_&]IaR;VO>c>5gU\^&f8BaYSaJL=EWe@UN>.BEQHWZ_
fY0ULX72)ET&3cIMB=b^@]K:RZ.=+g3HO2^;B_Ua2[L.1A,\&)0,IbgF\69#[R;[
,c#;)KW#b6REFMcYADcR_SLDBZ,ISVDGeC\N1YU#RM;=eb)/Q>cZ]H,TR7F#M:_8
eT5@8MF?+7W@2Gd+:T=I@](KK:LMbW+Og,]d+>cZe;FGJ04V>9+1KM6,<T-I6)WP
/)X&&ed5P9[f#OE/1ON53>3&7.,OV_]:6PDH<:)]M(I&Jf.4QK20#?B;fBQ9:IN8
?5TOJ/.<<4_5DaV<PQ6)^g^:\ZG;Q&[Ag(MfYUL[]6=.68B[7Yb0EeMN_a0eR^FY
_J:;_;GK]3ZOMV9Z)4C<L@65R]1STeFI4XI12O)E;00ZO3.6K(?5,@?OE#f8,D^W
@bb8UBN(ESGdB]:14PB)&Jf3DME7&fLYU&4](e1J,M>4H92>_C+I5JD.\8a0A?)K
[<T1DN==<62Va=48ENNR9<HKO=NB8Pf1CFYYaA1VBFcL.cFa+(\3[e\Ib9eYJM^^
)\9BJ22P,\5[83::[,cTCP(^O:\)TE,/?ec.515+;8W49Z-/N?=N7?)[7S,DYSL:
\.HbaJP<Q8Jb[8/HE63V):&._ePA;#d<W^A#QZTRY6;:]+C29NUFK-_JB-_[FX;.
#?XNPW8>V/g,PIc6,5Sa@3_?9ZA_VgX+W93.6a4^Y-#8;8Q@dU[V9Bd)/8)[2/^G
Z\;@c4GY]d8P2JS8M6&M8.M?])C7d/)BBQARUQ<RY2A_@TNS[Q2^5JM,K3;:bf[E
1;(+1E;\]6J4)T);)W-[fgR7+H#DGATVS_#F>(3VaZEX&<4I6/M;cWfd:NI.89Je
?2KPT9I;1@82_aZ02(ZDR/9HM4GE[1-(L56]-N7d=g,P172gJR2f5/R?8#)X=d[1
,L>bGRa+//1[O)=1H?6[J>fI?Zd3CcS^#;Fc;5\d/4b=KEK@ECAIFTU/+dDLCKB9
:VA]_a/8a=K>D47PA)dEdLbJ<])J]=HNNf+I#:\?<X\eGc\/O)A1D]1IYM3IDC=]
FMY\@BGAUL/YMdSA4KMAX.PZZ;Yc=]6M2@QTWf\MWc#O(?MaY&JB3C8DOI87c=V^
-FETL+F-aCTD1=8W@31?dYaPXX-2:-Hd/SBT:RN4?NaaG/&eF[dQZM#86YP5W@6N
2V;dG^FCc(d9\T?5_aUQT.I.>]bB,TMH1NJAV)eXA)LYdY.BdB)O(2H1^ZR;ZcDV
W-<I4)6P9>4PUF+ZefHLB?X36Y6IXOaefU\4=6N@W>T3gK;[THZV:5VgIU_GT&OB
TdYT&[?(.@7X4\J0L:gZ3MU@)Y3R7g,8DJOO7R]ZF:1E^XbA.fZ_=A]\.Z3-]H@M
G#IXVML?TcOeHMKAQSX;=,EX=3[A+(E@6M8d.<N2P8[F^Z4&ONH^C_:K1QcO6#Ld
O86#N^0.)ISZS5\.@fSVXcZgXPBdMMcJeZ<I\4#EA:X93(RKA?cTd;Q.KT@VD6b,
I<U<//_d(B&aGFZI.0fedgf6;Z1Kf&CQ=<&LOLBH(PK\+\.+QLG((>ZIfaKC>;(g
E#]=#3Ib./2G)S5V]=3U\(W@IH\F3K.YAf87KGS>DSC/?g\d-0e2)XM9(gDEHYe-
N0\=HF6Dd4Aa>N1\F2fEY0,BRL6>Sd^PeE>QQ.QZ#NSBB+S-48B3)EffWA),2cXe
NZ65Ae#T5RG[f^6N4DK_V8ICJR3HVKaNWNS>@3aR9dG6;CFID9JY6E>(XKa9-7aN
:1Dge@0d>VZZ2H6,AGYe9G]Jb7RR1W,7B)9)cV9PX47(KH7&W6Z[OVZC\G9>e(^_
J6#3FN17-Cd:P#LH:4?5:PR32(.cVO8]R8\U0I_L,]gZ5E.dPB^:eB7GNZC7gT[(
;8);(ULEg#ZED)-/]YQNM=/,:>T(\8F58;KR_Y@@Hb3<@(:7:>06ZP\RWVQPTXLI
5H^/_\\Q&)P+79QdTX&\d96.0eHC2&J)>.TEA]/CNg?S;(O4dH6Zc/aU4gKLLcAY
M,?])UXY.:@U)K;@BJ\^U?UB(M;C(R.)KY8g]g2EGa#U5,HRB]OW#U1[@/Y@#_G6
NAf7&QQ:@D17-P;Hg4F&<H(g,:LSO&NHgc<B3SIE5WAb,7E;1g3Rf&,2Y/5ECZV.
FUM0&eIBe#8.f-Q4F5\+C2d38B48>Z&>;8U)A,VFDN02&K-21><_N)>BYeTT#X[Y
B)H5Nf<,1;[4[P@\_<+5N)+OGQL3Z_H+9J&3CQd;c85KDJO,7ML]]?R=T0^:F8ZU
\@P:E0D/70NEL<?Z^GD2/;f=?6,cV^BMG\6aS8Z4WC\H<<0<U.]I,PE@VIUHUB13
+@\0TI,YNMQg-&-eSFg;7[\3E/4ZIBAT72,C0:b-S.>f/^cKcHgVgDaP4P69&<TB
/V]FBH9X^,Q9^RaPK]>?SM\b)H;c,--.]0.dD^fD2Ye-7I]Z?5PX,<2@:0AW@B>4
884)gd[@>O8:KU]dNCOI\IL:#-WLYSMIG;4>_,9OPEdNAQ/^V1/R)M-LR-]H+(\C
cP+R/<OLK9R5a>\d0F-NMEfGVCb4fS_bU1]97JR;,W1\gZ6=cB#K<GL_G,QV5/3Y
R.(_,,>?9(C.d9ZfT0aGO;)OC?3WV)5Q^.3dJJ5YA3f^<A:Z10&-AI?Eb79/FUS<
B[XDH+8RE7.4R.Bf[_&<014Nc2XW(_6#OHWR/O0ZB;II9YC0(,?bRB87M]0(1U[9
e1NHAWTbc5]@e,fb^IOc+H/@dI,Nc5.g:[HBN-XdBd_CC0fH^-NCbKC#RE_>,]DQ
E4+;f1OaP27.e^.CAa+1-(=AJ7<4]be[RC+5?F3.9HVOO-V<E.4bI;P2(O#:^YBD
d(IAAS-#I^YX^Y_)-@:]9D>.dN_cW^>^d&d?6A[,^#&#:U(f7TO#R2beISge&cM\
:?f/3&O&&_C,\]cWg0]/0S.J19P.UcgeR^O+?V#Q,If^8.6GGdFA9BaUZ@\P/SE4
K9NCB=B&KDFb+ZgH:/[43#UPOIaRL+a+0Bg(R3\:K[ZZFB09I@ZZUC3f[g1V19?B
S8LN_TW=(:>_@&7O[[?4.&H\POc,bWCP175bAX:Rc=BcXLPX7>I[4.<aS3NP/0KU
T[De7Z0:YAO7/8&MaBY^3.b&-7KOE1)a/_@HX(&7,K4=U=FSX+E18EINV(TcQB20
Y(L/P@J?I?X=9aIJ<HTHg=RQ,Q=6/]XM-Ad09R3>.OHP#K3=b0:D1R;A&R-eMc</
e13f.3GGZOE<194D;XI?A?YN[Fg0K/c1PcJ>ZNb(MJK(]K>W7REYfDD/U=@&5bH)
,:baCOeL7FU?-c70_Z\)df4.)[B1WUWg41E#D\fLUcIZX7Tb-5[-)V^-)9fKYN4G
&KJ.V3(J;V6Y-72]UHL0FBA)IM&\5SY;1BHS/:2;M;f^FSEUF+K.T3Qe>eW:JWSb
YB)#=IU9cWIbHdR/VPggc>)D[Rf0U,:U8P,[#&^I1QDHbYE[8KQ(_8.@P&_+XO56
(E3)7?@PSV?b,1/J\#B[:fR8\WYc1O-Y2QE0^.Q+F4#24(3J:<GBYDME9?@fGGYG
LGcBPf,CX\JA?<I6L<B,_RBTI]Zd>9M,VNB\d9fT7eMaP0Y):XY9G^QTWZ:E3c:O
JE:DU3;/_g;DD;Y.F1#[Lc;P&E,&;dDfJO((a679=&6eIXMET,2D=H>K@DH)0\R(
<&=.c4LgAeI3[C5Kf\.NUX0P@ePSZ0/9<@JJ]Z+5IHf6YHF-@?BPL=Za(@N<QJGQ
\BAUZS:.38+WM1-89M@5#DK+UPeBY^?[:.d>5TIBd:@.1^<^5a;0+_cA5#O+Q4+/
3KR6)]0OWN;UUI[;e_]aTDSCLB3RP\8G_Scb:Vg=/d60+.c]H.HD#/5/J9Ta^5MX
)#JLE]J^H-TKM]ScKaU:5G,58/3Z++IE+6FUHS?+061UAf9+]dF&+SFe=HT92f[#
//)OKKS,-00NCa<49@)bR;XQXa&@;Rde&WKLg?757:E-(2(3TbQeQ.1b(K#Eg@/O
&5D]9;?OV:a?F1Vgb65VZ@S?H)<c?>@c,\?S[KLOYV#77.c<ZPP5:B_aL(3\fLG@
B#ISB_R:1KH#GH[S6@E?\TP]2.J(S_DM+R/WeSF#B(g>NR?,E@6gO])?c,[b&Na3
XR@M[R5<V10f<4XJQa)CZK)PX_)K57_WgBV<3T=C)<K=#+9XFNb,b^4HGTUQf039
]G7KV?2=X.WERO]1-IGbg,<MSUVg/T^8<A9bQ3&ZS:-#>X<R&4L>Y8L0ZL9g&JS^
EcL>3/Ag;9<[=7A-QK,b[bJ?OZG9JId)B^3gcbb]4f=BN)?:G&H)Pf]NR]fAZ4/+
HP0O)GK=[g7;R<c^Pd/T)g1[\BH?2aK;+I3/]+BdN^J^QI,b8U\9S[98RC\),?[_
UYe7Fa&[J],_;bee=MgQVY;:;SE,9f^/>YYg>4VT;^8A6^f[A;#(,2EI0RNQNQXV
&67fddXN?0V1RY(/;cKS;V=deUQBSW:&>V8O1&DDGI95FM37dG5cRF/5M6FA3R6G
^O#EHD;g^#^H3812FP(E&eg5V#:/RVG.e._H\UUc,>Wa-=JM_dSMDOZQTIJ;b\<\
^8-FO;c[\MB3Tb&5gTRL/7c,)O;UN]a)7Q)IKPRAJJPB:C+-&DNH^JKTDHTB?F(#
&B0OfS/EJ>XBHQCE]a._0cYUZb8ODW1IMJ\a6Q[Z@M0-;M&P7X:.fNf.(AbAfZP/
2LQJN)/[a\]-&?7T\5E&.ND5V[:]5)2GBbW]#-ba>V,O(XOGTI=PgR4R.FK>ZR-#
OWXWJ3V3I-]&]b^C?C/gE671W=Ec#K0=dYeN8QP0F..I>XU,>4dA/L^8c;OMR[J2
9R(V&N&gJK+=8(.)X=A/VSI5LF-.Ec[S>U@V:WVQN92E):(ABCGXK)ICHf8;#2&)
K\OAC?^=/S&XF].a>I.R[KV;4K/425U<fb9B&QG[bX6)(N31[T5)->6,dJgWGV1[
8aV&S52^\dSB8\V<2]4bb3+D2JC\)D^SS4=^Q]141L,)/NKN0C@#G--,)dY\,,1C
V7@_[a&JFf(#;<BN>eRKDae>:_C:2EHED,]C,]:ZT&-aBA3C1Kg?3-b@Y</F08\f
T)VW3/L.J^G]POa;_)]-:b@Yc?+GIgfRCH-EBBg[-S[Le>4g2+1Q:NE,C4B8d26L
FCYg,7I?SBAU/>?M4Q0)8;[0PV=I?OcW9SFNKTPB4XPJHPDJ0b6CUO[:@NT()C[[
I#JK>bW)J2e.4T\8eQ6\\R+;Y+6T(,SYEWfCBMOXa(7M+L.,MT8VBX9O,N3PXg:E
<.AV3TeC,EDP\fZ,&M+-MRdX4#(P,6MV::e+=PP4GNKK.d<NeAR#fI9]2;^&V1,O
@E\W^U@RAD2c<)Gf(UXS&JM4I6GULceOQ^1D4G1J/Y?CBH57PeHWdKAd_2b7[=R<
FSWWeBT1#;=\J2:PO])^W>R-W2g-^C#-[0H-W6CVb=H>2KPQFSCI;I<1/F(MO5O\
ZXY\/U:HAPJ,C[A]9LA>UXJ@SGA)+.@Xe?5I9^G_5;d2L8-CRL^X^LV[M17d]V^b
c4VG.BCH71HcI;<DIgc4_E\3)IBYDJ0=ON&=8\>;.L6HV_fdY2Uc1:<:de9Y>T+=
NIL;;GPIE,5)B&P<)eV_H&:WIN[7Y3E]BUXg7FAPQ>cUY=&XGPYRYHG5DbD/9D?b
YQdI1DYeSV^bLGRN,@++R49I+3MC3Eec\^JW(9]V7eb#Y^>U#d_@]J[MU74152>I
X/?Va,?KJM9g_dg4<SZ.,cVB,GE[I\@?:.b2M(a_Mb=^UIc.7_,DR@0>T2RUGB^N
1,FF=;YfFaDP_\FL6^U<8XA#ORR.)CfY5F80&J7PJC\K6-.(ONe63#EN<;Fe5Bc(
YR_.-5eE#,c#Q5;I@NF3c@WR\P1cV;H^faJ;MdBIG]6+FMX:P9Ycb9L1<Yb/K1fQ
09XP6g8/BF#0N)\=OeE=<.;U]PL.<R&W0aBFObFXA657PT;bXH3(/<9SYPY23XYV
f0=8R(&I[6a&AMW6>/[T+aK[W_c733(Sd>IS00CFMPJ(#G)5;YHL>@H9fU0QDP./
cbAb,-J?QR-aA?@Z9\,0g=S)^[Xd73W,E>f/J)9DG:5?1(bJ414^W-6=b/LJ)>]d
(WKIVR?-gF,7^--X@_92g6/G9U(JXag&5EeM74WV@6SW7[d@1YG[;+\,ZHN,[V,c
@R8/Q1bVCf^2/HJD:WJW,g<[O?AT11^)UWG256FP><4d]@12I(Y[)DGM@<c=>OP3
;RHgaZ8#M6.75^YaE37SHeFG<c_Oe&B6L7OGR\aT#XD&;VDY\53XEK9fAFD<g?<I
0SdX45WF)O:6?9a>CgIQQ23bR(>6T)/POTYgG8>.)B[)YO&6e0/4)(9N,9C)Q2+=
P;A?R]b7XJ5D^1F&<P[EV[+[:9bF#5E[XUE4(f3B&W8MM.>[IV1aFDga]@M9W_WD
)Z]O^gEBf@KgDf4CX6&d+SFb0>XSXNZ,XT1E1B.4YU/49K;5[,a(a77Y\PPY2P\H
CZVWYND>SR+[<HRTRQLcS9?>N.NT2&dag6;PMf^a8IB#d2BSS+KbC)8g\N,Y465e
a)<M)bJVM/AK([acG&I9D:\I+>S-4T>??T]092Y&.0Y^-1ESEH8U[_7V<N\dI<A>
VKC7UYP@fFC.:a/C\@UeII02A.a0Q:)5IAP14)0GX5aN8^7)=R-DX6FX8bE_8@=I
)b>L<a,IeHL^4C+@Q]8[@:/W?04>.I1ZTGR9(OYVI8.Gf>b#\<VfSV\1BMfWd0_2
Y]dEfa;P/&AdgU&6d></G9H(ZRL/_E>\a>7dN46f47<,fTMSUVD#S?^)S,.:OQA1
C66#=DJ-Y2Za7bXf@5JL(Q(I[I58;Q([ZfP2[c:B-MP9J38L7KD3a)#;X<PL)XRa
6V3>M@d26\IYbZBP@/?C52L.UH#;>XW+3[J@1V?KE</UM(dPfF3,f(R\80\T)#?@
\RUICR^a#S_d/A(;RH_KJMO<Yb3(CKJ1QPB+\NN7TYPg]Lg=@QFee-6(H739M;H4
.;.OPFg4(X#4HdJbTgLQ8[0Gg]]:7FWLPT+gCGbE?0ccP;2:(^N]7E:V-Og3]=/?
gX;X;6,_E<.4;#-CDBgT1EY@Sg3.\1&c8G7gdT+Ta=+JXXT_[(^E<1Y-,6;R,Yb3
W:PC=>:;<9.f<6PJT+L640L4e>gQ=\,eTE\1+.J3c^]O[V+L&3M5.BIQe1X[fXV.
/?Q\#NVJIfG-=+L3f((U<:YCcMNH+,]:_b60UI<OTU(_3@CZ8bc_]@6E)7d1NCD&
=aI;4dL8ZN2N:=6@f,]85/_^f5^:;U.af/:3AO&?^a+G:K0.^H&5DMJ8S6>ED37,
T/[[OF2V1DC&<)@_5])B#IMC\+9D1CeRTf4AU@[G[CCE9PCXg#>NOBRf0DgM+A6C
[HYP;fK&V:H4\-e@VDSe,O-@(/Cb,<9MLCGE6Lg_#A@HgBIScXK/Z\R=DDV6Q^D>
X8@70W9QEFe[gDV2ac+;A/c67NYc2WP2^K#=M?6RVeRU\=C1^6(/Qg3cUb5;?6EF
+)YD2P,SFOC.aPS8M7[S12-aK?]Jb7?gW:5cA+#1+dNKd1+M)/&#,W]W\4TA@JgO
d\),f/E-b<6CKM7L3O(f[&AJ:K-2227K4>bR=L.46eHaNd1I;HE^OUbJKXM&\V7S
X==]<-7;Q:KLY25:W.J(cKV82)PCG?]/;fWcW1O@,gGO6VIcBULWa/[NME;LW3C<
cDXc#1&UB:DgL,cbcI@WcAV#PeRG2HK4/9gbR8<YGOMWS,9+4EYPW<7944LU&J:b
MB/255Z>ZZ^PgD8NbbGd=;D+a9,XXD4AM31+<Gf=,G46)KM./0(gbM2+R2,2L0IU
=,TP?AR4/..;f,f<d>OHdCC7[JM-&X-]2NR2_&X@/9PU:SM]B,:6/(75W4EbI4?+
.c+Yc06gTUBdc>OP.PFd=bJPJ)d:RgJ\F:/6Y2X[EV87?GMHLHB[cfNWf;Y<<+ge
^RMN:_Y?M+=4Z&S4(N]EDfSE_N=3-4QN0QG39+g&1d/@Y)J88WA.&R#,7LX^BLL=
D[4d1TaU?G7a+;0eL,B=QZ2X4&)QDQ6g:Fb-]g,.PB)U-X0f;AB\?;cKKF]-CK/A
20e>IM0Z&gFHca68)d7Hbb-=/UE;V(_MCbK2)@:D-df9GUebI?5M\5XNPA&M)RGI
Y2]b+CeL\TP/L7QDK306XU(E8.V-T1ZFL:-5\Z)JAS]>5MEN5I[ZaBBU(Wgf)f\B
>N#@I=^RQ,dVK4X:V6EH_RYYXR3.G#C0_VR(JBg(AV&gfS@^;Y.PMPE2c#(8V)cO
ZZ=SA_A,TC_aJ??>>VH8Y055.?I[VEG7US^4E79,86+MF,1#K.9XW,e)\,TYcLCC
7W4TF]=LUgVPZM<]=VL:SZTPB_SR]gL&]T?<aO5JVec=W5RPWcN^2IO,RJ0eTM@C
df3@6DU[f9,(-NY,6OW,.M?]adH>DIRS0M_<ZLE0;XF;:e:^UT2KBReaHP+R)H\F
7GAY(<8S,<@L]8B\5I&)X)2X;eIB6L,_D-IL9,bH<NK7YO,U9^Z4.GTg5PL>,@?H
@4M];e(6fW[<VPS9IQ3+@UQ<&0WcB[PSQC;g+OJd7P]AJ,^feSF:e>MO[YH5KF?D
S6V#aVBgJ.L[aA+7(fNECbagBSC;:>b5R#V:gU5[)/8KJLaYN<7Lf2#2(KC;dY-L
Ja93)VMF:[GMXU2MIBa74_.6L;MO3/:CSMffBbdH.,1>(I1G/\,6>g[09&(K4(d-
KB+GaN169VJ+c]aG07-X]F@O0;GTXUSee<HYU@R92N:S<N;N4e&WL[NPWC-(F._c
5aR-KKT8Q#d[f?Og8\;-?<fO&#;e@OSY7)f=,2>\.VCdOV4]K_.WQYK&B&)BeV-.
\>ef[f>=fGgQba?dDG0P_J,dRfN\)1NeN\XG;,SD.7dP&5F(<13@/6#I>N>J,E9(
WNM[QY,fU]:LS1GMV43@+_]EK20e0U72>1<b2NY,Ga4GK1I1J0H\g&-I#8d@D&0\
N>EWR]VbX9T)]UY(J6L-5>:1?_)NaJgTRMC^E5\4K+VW<<9XSRG>SFJ+Wff6(X1V
DS6-=_&6e(PG8Z0.D+EAD;3BUV_8D<4BAgVDYObJ\#G1NQ8>LC(A<0P&gWLQfK6V
E<?Z11M:>f>>B?43P[:]R119?bVXGXL?9g2231\Y>&YIPR/,?6g<3Gf=QfEBJeJP
OI1V_0f+;=1ec_0_fK=/&UTGM?=.0KHLCC_XV[M3SC@>2@H#C=KCHTD#IYK\gLRH
\Q:5-0JR=)DWF\E+>_>L<KDd67.d7A/LQEZSQ=6@a(<F0KU/2>UQQZ&QcE(fY:GE
:bMf-D>KLg//+\<&S5^_R&@8&J6ILZIGT[:fBO8RJ7Y-,a831>b#[8,:OX4Y:>2A
_LN]aPNHCV?]D#]=fS&[ffI;T5beWUU5AZ.^CP0B2e;K19[06Yf_<DM_3OAC]?W1
B:Z?8-XYRH-0CC^0;&.PcWULC42<,##SK&OSLJD5=O/M(-GdX?Td/L,f8/H;#)GL
>8HbPV@3-OWaNZ0OTYFf\]H<7Z4TQ+38YW3g)eDF)#O\M/7d]._+-PZ(RN8cV5YV
&>E;&&N^P4WQMSU/S[_A1HB8NDJ6<MSHJKIO\-\UXcNJ(/b1DR>QgK[7\>;7PR],
GZ]1,IYO9bC8(U#f:X-)URIYN+(eL7d4ee:8ADI&GBAfBB6W>D,Y,3?MO1Z@a5\7
RHHD(&HNNYNVNc0;^]T6J1XKKbNTE=M/]].c/P^JdH5)1[]>LQ7.@f2B/2R+37aL
Uf^A3.)_b303?2K<8&-\+6^)<f@DaS4N->ZC/&,UQ8P)DEVF)BWIK;RgM:Z>_bb-
673\Fg7GOLXCbUIa+&@(+JE_TC@(;<U;Kg7FXYgVcMEV946OBRFc66R;V2=a7)+)
4DZU\\BE2?f/N<-RWU<E;W#Z/SMef4Q2A8/Y^SF+bB4RB06&\)c@1UU1\S;,Q&]@
3OK0,_2M#/-?NHKfa5-=8B#9eT54/^Sb36@LYcd;=ECQ#Y(&Y/LFcDC;DAO24EN&
UWWQ<gJR0SW31[]Je8W;eNLS1VFA;:.,03fL6XDVda4C^+<YWXWeC@YFE-<bV=Q7
ECc.W@e4#7JUW#^R_SD4W?4ZUK=F8QRa8DD)DCO\Cb&T.DfH9cgTR#>-E;-<?5X@
L2G7<Z_M2H7^,d2G9:H8?)([g5^44K.OKDP#ZAg/[BaL,Md?a/13_5-<NJ=(J/@I
>3,:?&&+K?M#J:Bc@IFS5KHVaLF.48?UZ]Me6><39Q,EC-9g[X2GS_383+1VJ#VM
A?^^3]@f10-aZH(+2.[-@D<MN\eG1-9;UN+=3-C2a[bLb/>,NYQ0LX2(H:M#W:cb
(E+f.G<C??M&P.=)QSFN=(9c0Z;S@L[M]d8XC=eILFG]Ea)AM)[4aL&3U/QUEM_g
I.AB?S,NK4AL\7Jdef:P-]-]dE&,E\6,c&db\V&CM08M<=A>:V5VUGeYc<F+LI3H
)--@9_I8M4V[CDXM+UfT20D3.?OYP#UB/+?]P8f;/\N>_J3#?\EdV]g+?cBELS,?
DfE(5F+P7-K];4&5[F=<TQ?81;=V[S98g-W\ZFN/D+K.6R(0XF:2P,f=^)#\aD_7
Q8NM6#H<aXU=eSD)H=IgNTI2d3d79?a:OJ/0LGZY\bI;-Bc#NN?fO5YLcIa6F8I@
]4eMc^;R1Xa<_)?A95?-OS&3U1YF6M>1\Z4H,)4^?cKVXRFLY/-:ELS3+6\];-PB
^fQdKOR2SRSFJaHZKRY:34\D.RE-;d:25T1UScAS::(BA,_Q)#>,1&>XI-CLG217
/>I]Ub4ZK+H3S?OR]b=903LP,&QM.K[F/Qf.e.Ze5ZHWK:2^2XH2]2-eCY>;\&9R
X(6-=IR#UGXCM[Sc;e[#,cAS@c0d7<[C1@6<78@gbYDR</0K2PIG.9dZ9HNYJF7:
b+L+&/MGX3S/=2=6JOg,e^WNK4ZEUfA?7Dc6E)UT@L#17<86ObA(b26AEZO1C/I>
eE_]TfYQT#+WOOMdbEJBJYUO7G0TX?UX77&71O2cdEcDVM#&W=2D<L[50O25Z,#_
N]fLH#5DTG8X<###&;_-NP>O)HA#>)g/=V/7aP4cfR#TfFgX[[d9V(IMaBWaTc.a
,gPS@-#BB]M8R-_I+XZP.M412J8\6:\YeE+d6[6:)>ZL92eR3g/=1BT)&D(Xa<7Q
5)af=D1)F.8567S6L)32I@Z]9cI1(g.14)A9M@Q;#K[Y#FD8:T:,G,[C&aX\D3Ce
^(ILX([MI#-a:1Fe]0YC\\DRbJU^K_+DBc]DQMGTDO<+9IJQE0#S.;+(.Ke,.Oc(
=@-_JXeQ2P617,CLe8gZ:/BSb&@2&_=^>B\J@De9D,VQ2?\CF[/O#:0N-NY\>O@_
HY/(dX.F;cS^=_SUf2@YD6B-XL<WU^UV<b:Yd6c(MRIJ8Y>QT5,44T@,5bb0SB>H
+Q&IZ5+U8a3]U&GCI0W590?&8>IdVMX0.J+,Y0Db?M9\D+T&,#P-PY4cf_Z#088Q
?P<6eBB70>;UJe.JDI7AJ<c#9ZL-1>-1,=d/GT58S@29G0X9(dU02)TagP6Y62WH
3K\A#Y89_A=W@>K\2f42c<[N(,\7P<aU@\4^2).&HeYJFNI5g7X&dX)8.:I]WGUL
#RM,S=IZ=b+\9TdV?5G6H.AXEOS7]a)2b=[(0?SeT92:)8fDI]?<@_d<F@(KAI2(
Y;BWb=DeJ?N.12Se^@Q^G0I=H:7/[/e,K/gd?Z5/ac/S^dN88W&e/NcNJ:Z6[^d>
]8^BLF9?(gJY0[A9[Z2T]/8b-d9;)B1SERUD)JM?L4TL,;@L<#K,APa4/d;P_F/S
AQ\(+aa-=@;96E1H2-A^,MdcZN>-#P6(S7D,T-0c@U<6LAQ+W]>:?/XBBX3&c.)?
.2NZS3gC0b4WN)JS_V3K5a)UN:Od/ZbH=aGEdZCJP#9;Ea=+c(d?3S=Qa(#2)8PZ
EGKDGM:\+=?UU4>KWM)\a:^^bUeU6G@Wff2:+8LH:ab@=POX<M^LZ#ZVN59e>:O1
W0UOMVAQAMKgaOJ:-#27:8+4M3eWXUK53F:3A<d)&=)3.b=LGD[<.Y;^F(LKV)FE
Fc=&;A<5R>RBQG&RYOH99US[X(ST:=8HP5>X#a]gS^DQ_1:<46(ZdJaKBVOPI^=P
;CbLdNLd#+HK^,bf\&^&AF503:02G/W+6X,RO44Rf=DX.B1?HFK2IN?0JafU0#-\
Q/c2[UO/\6d>(DDAP>c[@=(3a;E,>L4;FSc-McN+-4SY[)&-\A8(S=MHE8WUHNd#
aX=[SA45HJ)F=XTO]XeR^d&X71950QMH5O?P)<DI.?;SJGMOL^UT;F1X1#b39b:f
9;fPeG:^5;5[J?CU3,XTK<L&1I+@f8?_^CFZ^=G8\LY[DbQ)6BA1fNP+5]^/-f0<
RO/eR.^aX2dRZSc-MGD\]KZ[VE\d>3<+,SRNJaS3f+,d;7SQ47(##bA2C/=D:#>I
/CSYXgXSc8ZWGe0ge&HaKEXO/f3\BcIWbcWW=,/2)BEZ=dI8K;7(U(L)cEO4SZPb
Z/3P,]D5FY5f(F-e\g8Z59Q(R#f#EOC/[>(&8J?Z7.;De5>WCQf8>9VN(VKDXa.N
7L:^M[6M<N9deX@KAOVe?C0>##9]OHb_[W/N/JK)Z99[KO7POQL\3e/P5(VTT8,@
0GN-c+N0W)<X\RbYYR]X:,&dZde4RDAF]0(-eJ+MVgTgZ)4.+OP=IJ0)>II[&a.#
TU6RDKbT=RKRff>a/?0_QWfM&dRCQWfK-?VP645L=4SYBfWOMYPOg;04QBd-[d8>
^O#M@XV\g29N\g2;7[Z8ET0afP4aIJ+[RSCH>T8+a:7BXRS7c&Nf[_F1E[dL/X<\
gg.IZ@G\I#Q(_fY^,bfI#70[F?U39G&\8[EEg@3]RXRK22fS3PGFP]^6=O3.\+;N
Y3.S3[ece8@)fMA<(1<cH(+Z0ZP6=L>_-=PP@X@.[V9=@]bdLUU-CKZI<<a;D\a:
gFOE4I\d\TJA83Z?Xg>5V.F8:^/(K]9-=>O2585NbF0X(0D[7A@9JZ<SG[/a;IFS
6F,fM+H;1>3?G3BO1,;/ZV:cRV]1)AE:J0(f5KFN1eN4H\@S1C0SYTI1TV>c^f2D
K3TPERTR7V#9[TQfNJ(WgM[W;FPR6LNYJVUULbZb0_35(Te]A73TMB_:+9EOFJc@
QJVL&2Q2/#9(X8ZG,@PaGaOfB+6TH]7E9+8TdK0GTIO^<5PaaVDBQX<T/2UX#a#0
CAZ.aX2\RY(#+g8FLY<<bbCb,7ON3>MDKEQCPFI[O<\_:.6UO,cI#4gd+XEUEON9
\J.4)U\IgM,#/(IR8O@eD=-XMX7-MRcX)>T_5J.D4#+Ea1bbcD9?b]Nfc3UTG[-4
EGEOU>/?)LE0aUKF;P]eO-IW4=S3;>E1.c=cWSD187Zd[I?&VGS^ZcG4D+K/LGLO
<NGe2Q5>J#f/Ve6_D(I9,65#OR@^?2D^G&D<T=0Q4U7dWgGb+O124<E?WIV@7c&9
&3ZU?X2cgZIc<-,[?3@UPV)F>8^1,f_a.U<3?b0TIEb_,MZNW&PHCAa@CR++<=9]
;8;EV\d-[@JVF^G+S@A>C0;U@;PH.LSLQ^g>2[0dQC<5LbY)AW[a)Nd<3J70X7cZ
Qfa+Q##&#C:3U.0LU&fHEBXTJFZBTf8P:C>6JX&/&R?(U8=;(S\P]e&W(B:UN0=Q
+P+[E4a9#F>5gM^,>RJ,IN5b4WY-ZS1AA<S,&=5_@e/8PgH]F8OD(-SJ@]VP/cVf
VNfVPUS7IZ68P^-#eDeK6OO3LGH5I=KC<7Dg<Y&gORH);-_QcT.[Xdb>R4TfVc=+
@dV\7#b4HF[J8><[T(;JX\7/EHc/YDD4_D;B/>J,F6=R;(^bFC]]UaaL8CZC1F(N
9;#a_?]N=3=gB/6OEP\U:(D17FY03[ffaS4KX();6P-A,EM#/SRJ.b&H(]J,g]d.
EZFL8e.Mb8cdKH9_a9Q:MWT.[R]<H59^L\C;(8(@4^.:Y[gT5Yc3e>@A?c:6AD?5
<0??&U-T#b&dQC@Y]?GY/]:e83YA35C<#3[F1\:TAbGFC9Z)f5ZF+=c1)/-(M99g
P+>?VP[)[DIdI@TE]H.d&+>8^;A>DELL--2:^cC23V8]&).-A?\NS_^IV:T:@e&:
S5Z.&1Y_-[U9[/A.HX[4I7A6K/)O94Gdcc#WBVb=<--f_=<^UFVZXfF7KI=Rc,OW
b(d7\67DE=dfRf[^@:)R3C>BPL^C/4&17f&MEdHG3N7cH?-C0g91,(PALg(665(-
\2(/WKB0M22b+E:_DHP0^=C+FJ_/#:cJ&28ZDL9=cGCS#e_A?C6&PF3]Eb5EVP?K
3^KA?LRMK\];6-P?#COT@(3=#Gf7N?[8\cNBD:0J2]4F#7+#-,^5VV62f#8c?SDH
-D>3SOYYEY5;O/[g&VC[51WE8HbCH\C4\;@UL_4f9?HLH9Y??g?YG[f@7-Q1JIR^
M;P[]7PeZ&,S=K/Z3J<<58O_.=a]6547UN?@VTL2(IMB([_>2S(O.f2M(0,<CC74
;-S7T92C/SVRa?Dc.[O4c<QT5W:F6_.cI7b:AUE)_^N.Q7>9(0=-dS&2T/@<(BF3
N59/9dK<?Be4-CU1[^.b[?I61/>LBYaYJM/bEdV3VB.BR6D762Y(3MZC<AfdC=dO
Ka:9?:g]bNPB@.DW(S>4V08U-&VYW2/9DOE]LYb]V7HRQ\_5V.cf/Q6SVAf7-TU1
/JU@)F>T_YHcX-9)\1S\(Zc[LV\8#6^0C9f1&JfgP.:&eg]/&d/g_3\gPJ>WGgT2
F@d>^HFd9U2/3/;bM^6S:TUN<C3<CG;IZ\C_@DK,:JgTHSNSb2H>3GA;C[-Ue.<W
BfHS))F8,#(Jg2&PVEKNIC8,9(.<Y1@[N(+^7P_FP<3HB[Q2Gd7QN;aBH(5NY2T)
R:,4(<DYRC,:Ee1fG]f[V3[&SdaCX^8>>Pc:R(e9G?JfV(Q=J,6_,]#a\c&BDdY&
Va;BeSZKLfZ7.D3?/<=@4:239Z]N<dYVa[8+MAX4X#HbN<BO/Q2XW9Y+#3KH=7fU
08^gHH8M2d30M1PS5:@N,g\TZ<^CDKYBOQEVYHTF>\YdKF=90-O8/MbVIWe[?c^_
RZY7>9.1S_eM7U.4@d<Y7P,(M6N#8\<:R\HS(#,bJad/)MRgRg88I_PY(9@fD7BE
J?ZZ(F9&.)9^_<LDV]>g=^Mb^HUEX&:ddG-;UC+2ffd[f^5.a@DaT]dV1c-=9^W6
>AZT[8;4DPIE0Q]dJDb):JX925\T<69E&=\^8eB^T;gW0O\KFX@0+_46/]b<.,J[
g07X^M@[3bIGL<0C_dELEHB=9.NHW?@7eIK#4dL5(F;QJ53)EPgN<#7LLECK)KH?
)IX+\34_eGJU7_D]Vd.TK3CKI:G6Vf_&3.(?eY\NR&U:^Z&a;N4-.0bK9-dW7VIb
EL[-8)6)EY+c=\@_3G2V6/EJG0Bc;/a]K)6_>g,:-ffX3#]L^63K3N#TTGQQa7KL
&_V4a@16((JUT9@ZcbQ67UMI=Tg50aO]4U:O^8TY<cPg9^cD\FU7?,K#/eX=3YHe
Q1PL)ZG0+LfMegb8C?AKg4QY0CQWSRY:)CWe2(:-&EC2&D/?\->Ja6D2T@MPg=/G
S)-@5.e>[PgN;.L]f[4AI-KV.BTTg<)JIX(A0f^\XV>8gZNTS[N2<&);@H>D\^\A
_R9HA3R)6D76Q=CZI<;e)QA&>+f23OW&&eA3OWJ,eIf.^,YA:-e:cG/R#N_YMMdV
E.a#<[[IPU,14_a4eU@N;aTHfC][/EgCJU>TY<(6PJ@4TJ.\YLJ&<T:@G:TdYK_b
7:bQ?_G\P9Qa:5gJB@<>60V?)E7c>bZL,Sd_=d44@aS)_=(;HJ&MOW32Z6X=:URf
CX3E1I(0HN/B,R\a+IDJGTO^/4?DaAdgRS_6OHfT)O0QMEXN.L:+;28[J&YWe/B?
/#fBCLDCQLV4NV>YHeM@:JI>eJ4TUeL#V,:&ZP>?eab)JGP4I05ZaKSZEA=(2:]&
YLA8^@YXR=\@O>E[GQ=5e2UFL=e(V-C):/PL12+\W9?76aa#8-WYgVD]H+QG\/T5
1#PO_ZaYN=SHGFM#I8?,JG;WEc((^e40U/P]^\>-5::(,FLR77SK0_DFc#VHgfO/
90U#>dX@[1&V[;&HN;?[cF[;XFg_e1?0Le2UTXgO_W@,cCfTJ^da4\K.Q.aCJ3DX
/9?D/@81;6,16C]-A[TXNVA+KFfb)__3^4Rb6<&9dLQc1e,&@[8B:M@S[2^e0Z@S
JPec0SYK,a@&_EJe&E:C0C1+2F3#IV&8aPG-4F_0_[Q[FY=_+a>:@eN>Cc_#aEb.
?f-DGc+,SR=.MNg#.,N3WJYNH]\#DB9(-)da_dKI<96?#U#O0UNa@7W9=S?DZ_.T
A9R?HMHD>(G.OE3+FR29\-370VI8/_3FX-(McA[HDGOR^8JD\^/O=:1)?/V2/&&b
7\Ba7Uf@.6(C1bG<b^S=U:9T3O,.RAY]@b,>dK2@4>:\+896NX\@5a?F<ETVR6XP
^=c9.RP:(36@>0S_2_TFXa<Bb3e<f.WM?<&_,U3+g6>?\__TIHVfIf8DM01,@IdR
f4aa::+LC<g&_FM(KAMU(5^BaQB7_7L6CeUN9MX.8F-V]^?2J:@+4O@P(VaN05V=
^5;OXC0]W:LfBRG._W7X9TRSCa=\R2R[A9]G,LO@fJf:V8)EKN?<De-YbE[223\/
O<cK[EEJ66:Z@U0JR#95b^4O<^Qe9N#AS@YULNM98S1,dL(<;DLNf0Wf6960O0JE
I7BRG3WA7P1+01S5f2^VdSWa]\QA2J<KA).HPA[?#._f&X5OC@=]QdMP89PYA\2\
&+>O<W-f))OYT9Q8Y)(UbV(EgSJ,]X2APOTd_2_&Y_,)]MdZIAC)3F7d#&@Ie=b6
)/]D#b.R[3(a\K.^2@5fSM@1EeZd.aYf3[feY/<7G:3AG<?B(ZOWJ1?KH94G^;7P
><g;a1^[,9[H/ZbXTd1#[X61WYFS:34KC;)H3cGM+8_6FXE1,8Pc)g<Z+/.<7,[8
O#(L<,+A,VJK_?>B-IXKKeGT?ZFI[0K<XIW8&2\/=7,]BGIH7VLJV#=&[ZZLcg1-
=HEY3YX#e@GWEc)L5M-SMV(PAFSaLg4?HGR>(:gbeM7_UY,=aX&W[H<Wde;Sd2cT
bA4MVDU3dAS=7JO4]-[.T[B7P4H_W]RQUV41)OO.QcYf\Z4gZCXQ-?_15D+\dNAO
K3)JXb_-#-Wc+>eL]P?@Y(5:cL-4<.cDHWbAWBB^&];?-g9G>Xd;#YaHBK[[KM^\
0G9U2X?M1;1ZB8VUdd9..&^deaB3,>a<a6ed&I8dIcfUSIS0bOWT>c3LE/8KCB3>
0bZ,4V;9Vb@c:K&fIFQJK,4&\9f?CX38TWN,O4)65fb07a#&NGL/YaW+2S16-[2S
.;^LF=2H.2OJ=@dJQbV7gCgF4H&dN-7PW2/F&0B+UFIg/VGZAOFV.KI=HIf#U;7Z
@KH7BK,Y(V3S:d472e94dBgeR8EVgGHE92:[EUBW;@?_Td\W@Oc@?/YRcbTS&DW,
MSVb,:-c8<-=4.X7GGd>>.38I8-RO7aeDCaUg[?<VXf#TFY)UDQ,.#C[_L.PK1E&
&0462>[@J(#JaCI;BaCFaIP:.3>P.=MH9&WRCe.fY)f,D)H[V8.?&e^--ege-G;U
?04ZF3A,;F8/d<ZQV<DfA6-JL<+;2T-DT2=1CTDNOaQ(^QHFgB)gFOeQf#IMAHHM
B[;&W,>fS;7X0<]Ef-QHR(9SeUCQOe3OM?I:?[/f-3g+O^0C5^@;PPceE.01I[OU
c>&Q&Q-4WMX6&H4FFPW+ZfR.2S3O.;9Q+E:C8PV6&K):?0=,Ae(]W0KgA:gb:KD1
MDUA-NPM^MR&.KHT@LME9[-eZ<SF/N+P#3O>Y,4&Gd7M1S:4eCcca.QL0LS,1HZV
)IgI+IgP)&^4K9,>Q@P+GbCS>/8(?SfgCW+RB5f9SAH1aR>SGgIZ@(dJK5(?8IP-
<&-,>.(ZNV4b8TH:JD(0^Q+/e](;KJU5N.,_C/0MLME]5WJ5A(8MCKeYcbNJ_eJ_
89TWZbKJJ^ROMQIAPLgeb6;..-B)#\;7LUf3CXf>>TX:8RVbRe9D,+(R)K9J;TCC
C-aTW,cETIeZ>;?NV=7D7ZD;XR(gQ^SQG#CCJ)8P>-Ed5_YKF]/BH6A4=+:4K2#0
>1VX06HTQ4WAOH.d5OF\Q.)<.YU1cLHHG,GcWDS:e1R_?_-6NBYaYTF70e1,BPA@
VJVZHBWZ=f6.9^Cbf-C11WR]f=S9Gb3aO]Xe0UZDYSE-68-gLWY?Gbe6a14,6WTW
Z_Bea&;T\,O9)fNc1SJ(ZTf&X:&bB#()gL@UM6^f/.^Ig?R.F<\,[NUH<(XQ]<0E
OQ2DDG3?-6W-aD96BWB5M\aI;PDf/e:_a;CBFJCYVb4ST:_+RJFe4YS,0HD&CCMN
7-e.O6)d>L39#F;;+ME9f]TMd2J.WW18^A<#O)Yf,\&I3U6^&_.e/SG<EL6+TM@b
]0?d>-E&VYM6>U:)MM^8@/YIbJc\3BBY4084K79Y31N/./;V3fFGAMLL2e70DRU0
42-N1#SA?g0aFXbTff(Kdc.c3T8gb7\9HMWe0A^ae:HC?<+@(Hge>/TP4J4@[(IH
8[IT_WO0&QSPYE)dPeWfL5eKd[C4Y0-0+P;F:0-^>+e5V^P)g<^9[8DLSVC/0b0@
XNc\BZJYZ/7B,^\QCcf0dWO]WB@=FXfZKdR1R)CG+OQIPC#f]bA;P697:;aAb+bK
]L);9A@REJ]a37594RJ4>M2)RXN#@JM>LRG=7&I3\>,@4;](]:JXRLT3?#f>?DEQ
0P:P9^3Pf_UM=5a;IBfYL&0NYLO:ONZG-PI;a8gec5]RE;5Sf-b+U?A4c25_=:&+
Uf?/KG4S>MESVAA^@P6T.R(G3K#egN\/6P,/e\gIJR:.AL-]IVfS1D\B:IcTM)3L
2g:DR]L+IH#PY5D+4W,Jf->.6^5b0X2P(a[(P-#5fNS[bIf]#()#6.WFW0d/YLUF
P^2./7BRGZ8O-_f_1=><2RaQ6<#XR;gGVM++&_[16cAcU@BMCXO3[8WZ2;PV<;g<
]>@fMR8egeL_?4E[7Zg8;39];ZV/XQ).L[7H2O&X<A0;I:;N(#>EbJIa1I,W0,@E
H:cP/8cE?RSdc4)b6)?HL(7A02H?=A<MWGM0-c))HbDP>03BQF[/c7ZS(X6Oa99W
IQN+OH0I=R6a+>R2R3G#751D1-X6Gf\dW;ME48S1)U2O7F9f#f4#&&b:WMA#F0fF
W\T0B5;Mb09?Y)5SN(K);PE75ac]Z5L@>.-7;1gN-Tc\17_72RG3SSJJNL3]_D]L
2,DL\LZTdN@Y1>UKG1V_-<OB:413;SD(GZeLC[X,VD;ePKTLYeBJ79)WC:J?W<60
88?1HPH:@@R.=F;=YgEGMEYcM/CO>8=d;6H.Ug=]P4.TLEU^702OL8-_UEPb#ZF:
7fK4a_A<:<<>S_)MNT<J7;<[DVf[@?gHC-2,a-)@;RH,]IR@e+(Sc34aHAaYZ0,Y
(]ZCaH?8.VR-bdWY.O^&c@d[NTI15DQ(5+;b3Y@e.)dFFcNO]^@2e^Yg-_+DbS?e
R+#+=ELdC9J&0)fU<5ID#6\V?+:1=c95^g3\=433eR9J[@;1?bSIW#+;L448KeCa
3EDAR9@E3;#HWFbKE2C.CL3#dI1FJWDST2A7a3Qe&?5SJ=O8.R/90D?c[;P<W4Jb
MRgO@:eY7B/Y_JO_&)40Qf05JN)J?78aKNJW:0N<Z=QbDZUP/Gd-(NR<+Za@V9?6
9&-(A8/YSA(b^&&YJ-@4D6R\P<dLRBY9_):F_UO5>YAYB8[cA)Wg3MW_P7OU+#Q.
V2Rdf/0a>9I,0Q.<P0a]+YH.BB2K.PU&6cA>C2fLJAg_3EU>COG]PA?&A>?&6Z?A
_J9a[PT1RU[\V5/XHB,16YU7)I?;/>:-XUICPFgBD@J]:-bI(NRGa++E#T4^Z7_P
&-&JBf0C3N-+SdHF(Z8;9DSD)2_CfG<RW@?7=H\68?ZSR>+9AVEV=STQW4:(R6WQ
Ce87ND_?R&_2(c;5<#AX55H:MAdO?X]a=\\(0>34VS5DV8UY0f23Z6BBe700QXf1
/:&M8Q]W#I?16MRTSdMZGge/A@_TB/2E)FJbEfC7S^D#4\#T[/#WE1Z+fC9YGN_H
a>EKPDO,]A<&MB[#7BJQR#WORBXCaN(GXe3V3Z?K(d.+gYFQ<ERM[(e6KFX#&fQ6
A<(/gD+9KK\YP3?,3?9L2WH[@205\:>L_Y?c=6dA+gcfU?&GD;(SNa1\I+<GI_\@
]#,L[d_C;eW/-Y-V\JJH4R0-bQ-J[DLKe9;=A3F0d:+BMQ-<E=TXBVY@Ja3g45Vf
20KI41]Jf(9dKM^NdOSVfN^LT-eH)_QRaWeURg(;eT-Y01M\T,D+<N9GZgHB7-E+
GO1#QSWFKI&Rc#ZCBZd_cX>?d_.DPT6B(IX2WfB;g<+,B;@a,S\X-YH]9JC=M^V,
^1:/5NMD[\>,K/T5\[7gU)<[eQJ?f9eNWg6g/_R8@)0RS<3AW6U9G>04:[\__A,]
MDe&==f.TQEJSf<PP/YdCWS&9\9G(4ADY(2]F-I)_RS-,dXXDc5;CK?FFK4NcWN3
V9DX9X8e[I4]EDNHO0?+Mb3])f8fDdX;a,Zg)^2TS8[JOWWW:DS;Vf+a(<7^]1_&
_W\A^RbB8W5L)=c:V0QHdF0AT]PQeXJ2R]JTd[&A.<1>>/3F(AV;]PZC=\8FM9B;
?JRT_5_7=_,Gd/>&)1=/SaY^;4>+O2\d]F5=?J)e)H;>7bPCJNV&c<96>;g@LHDW
b32bbTN,?c]C@>P]8>.M3;c1OW1<VDYbF7D)A3db[9G[V2.DARXG]#U6)A?VMT<a
RZ_PBf.&R9=)\TR_RDfRI+(7;,a&LTM@PD&/?7b8Ke,>a;1c2_FK>O(H.(6f&,Na
]_bWEg1ab#HT^\dUfJ9aN<0DH4HOMaU(O\IA?e3#)9+2;WM]FfMG&B\^W2RAQg0J
_LD3>ZcXeV]-6W5[77N2D?@33_@8(K0DfC@[42^1bLU]IXDHYA9@&QA0NYKBb8,4
_c5-E405HZL5.TQ,\I=DXX1.4A-_c4#O7@J1aPP/=e=8G&,,G,_MDI4OO3XEAW3Z
P-Cc2G+3T+W[WZSa.W#@.agM#BI]7Y-I-d_Z=J+SaD0K7AE_6L&W.2&5]b=@#M+;
P_Y=PP3QJB;+(5->9]e58GCaJ7ZX_+\(NIL[XNeN-Yc#>9E\?:5L;aS+1(A/==ZB
67=f1X@6.+1&XBR>&AP_55G:I1[e.LNQ<4;DcKVWA&<J8^M(;(KQZXMA7cB#5Fe7
B\U:abCQT9b/fM,e,THNMB5U+H66?RVOfUK+a^J:@?4XO\b5IHW2Q4O^,@ge@LL3
/8/&b@&@+4R(2W.#C=,Q)aYV0OFAKfY-;R^e6Vf#Z\UfXV4>7]gX8R0dU?<+bQ80
5:,c/HX.Y=Sf&\7S,4g7@.J)\(V;GS6R:(_^Lf]-JN+HdWO=a1PC_L>c2(H0>XV_
eL19VBJ2NRHF1A(K7>5gAT.FU=9Q25eB2V2_<W.Z>f3BN)OV^c,CXS,a]ZU[V=\D
A^@,)0VB/U9:EBUKJ+.?,O@E@P@.([aC-b/MU@ea7;ZL6<ICOBQ4)F&E<DAA-;\K
-@+8#&Y8EQC>f&e^VXF+-K</Y.b;S5<Ta;K(ZbP#/aAB4AGaCga:?AO\aR[AXd/5
=1T@0L\^]UCTaLRFODObQO-=\VU]+dB,88HF,^+030W=P)AO\G<(#F/OVgG/@++\
\A7(LLf,eNT)AURBR3-+e>Q=99B=^ZSLdTFS^(^&5=?c;cP@4@112NME(1cdaSQ8
eWHK3W?NEO]Ke?:3Y,7H#7d<2U1HMV--Ga/W:Re+5Q)J0HMWUEa82T5E]KMFAf@a
<YI)gC8aOF6C#];H(A<ZVK3R@>W5(L6E?/a01XT)D=0TVVU+V8IM-2R^))-.fZ0T
NEZ;T0ZU^^JH\>62>5de\/Q:XZ<ed#\b)W\\7CLa]8&\0Q##gDd960UB2B\7F4P6
?B=Z8S3B-Rd?3bR[L2YO8Ad01c+(<V)P5]>(@-R:.J+Rcg-R=BR[K+JS5Sa]/If9
YabEK-dXD<Ib\;N@U-?E-P_VZQ&=#>Z@[O:K2-d5@/S4AgWf-8-LEe,[<XY7OS[6
)Te)_H(T/&<).7IcD(aJ>8Z9]T.&Bd.C7D0aIBbMW,]Z^.gDVN5\)dJZe]FW1gJ0
VF.=+)Z1GPJMY48,83A;>_WD9Z?Vc/9UOS0J^Mac\?3+7geOS9HXTZ<8(U\O..[<
gaM:M1bC4\.CR8-?49U.RH#_TAg+R=FJ<^_d22FDWGM8.b[U7L@[1F?-E4g83Y53
b&ZGK=8gC?EB4K-Fa1ggLE;3b],eUDCDATb+I5GCFLf+I0=ZUO8KH9CYG5IEY;Y5
;G[-[9XAZ[RH-]#,\[+f0]Zb6G[WB>RYMdQLCa#c._)0WeS(?IV;U+48^FP.-V=-
1/g_QbU2=fFfe&Z\Qf,X0GCdIVP/UKY&)ST?0]GA_S)Ba57+f-BB7C)1EO8+S(eA
7fOIgg+>3NQUO.E_U7M=:Z[-&6L3#I&V(NgW_g:V_LKZYd8Wd)V6;WYUR@L4Q5)^
,5Td?g,GF]@?5CJE#<\#<6HH^WD:c7)C-e1&EYH]DT9\IFR<f[4S[aN6M98_QR?D
T-LcJA8VT1-<A.?8bHRfC_R^S]8F9O4>#)4Y+F0>MVP4D&Y[6<eD8A#;A:N7;TG4
MJ<2)a\=b?(SaG3)NKgT-A@&9JV[S4Z^-,+Xf3Rb(E;ALST/02^P^aR7=e?@WQ):
>DDI,M#TLF,C_eMP^ELR\S<CXe5cHS5A7I3T#H#1G_Mf0[,#e^AEc.,5DaFI\]J<
,GN]^YDg=#/,_N,??Q)bcCa:I;SG102=_:HUYY<]G4W]WL5Y<DAF7Q1/D-dM];E8
5?06U2H^1)AgT-a-FgYa^TBD&Sg3[7N8LJ+:2^f,XKbJC/]G>OO-I(7Ua(de2YKA
Y[cS-MFHMObCXI3<D72(FFIEM0/c3&g@SBADA;)\@&<U<a=H(6e[/+:/F^H)7dWI
8V2-(-\5g#e:ZX4FNeb:1N;+NQ5bQ\NOb](7:06>5;7ZAJ?>e5_bC+EFOHW-FK5/
R60\ISc)Z,[bW_8#A70aFHE\XA#H]e:EO.S4J(JXB^)_dHW-6&gTT798I.3(db+]
1bL\INBCBO+d:A]3VdR;3ZBEJ,gf]&AY.3N/Vg^MGff\2ELebX5)0TB><T?@Yd>2
8Y1W79a+C,O\JF7<74cC[.G0a@>/9J]>^_-.[B7T0/-AT2;OW0b2^T?KF,gQ#,JK
4/7<EfbS4KW:X]WPgIC]=MS)NHEAY<\+]?;VSP/9V5+(#09DHF8(Me_N.0+[e;Z4
DfHW4-=NB4ABLK_QSg+M/g6-1R?+<9KdeN:(+GF<_JF<fd7.?_;8GOXCe+a>7<MC
8\2AFH@V/<EZ\7&(K59B3;]DCF?)9B^MeLRb=(ZJKQ00<Ja8<?=#&dFBgVcQ\SDT
2&/L#]5ZZTg.dAPRca&<K3</Z@=>4DaXNWb]C,)0Xc0#I=bM0U5B@6>HC6U:S:&I
+/NP.WGPXN_W)54/-^:@fcc:a5gRIJNU+7I;]Yf_\1?EaGNT[_QORe[@QB^FB&ED
c>0_LgG5GC2<>,95C/0R&93ZBB43-F)gH<KKV5I6,SO:04.FH;A?45,M)dd:V+^I
a>QQF3Bg,PE)[Q)HYT3::T+/&PLQ(Q&.eSH0cW]\?c0+&9GaYd\^^6^/8DIXQS6>
)=:2g-E]RfMV2Y&L8\4,-.E<W(6Dd;\19C0A\71<e,_7d#bFB;_@AP6RWRF0<-c>
1BZgTD_5TFUQL4>VBZRE7\;7Zf@b;8bIH0-ZY0BZW^;M(A;D=HZ:?DX+8;X#(5I;
<b?8<F8a9(H<6&E],C/.bM8/M0]FJQF]R>aN_E1;O&Kf1^IXUR(^TG+):#?R#YZR
Y@X<9(AT5>NEIS7T8(4[ISGNY0R0O>;>51H2d,+4,1Xd=c^]Pg9;(==_G-ESfVI9
^L+C0V.((>:)UR)/^K(^@5>)MY/F^+#=>6A.EB6+G6aaDL8<27a@;Q,5+Q#UO;[0
,1^0.K6:1&gZ_HWY3Z[[/Ge[MJ82VI?g^^=#;DOJTHW_MZ57_[21.(,3=/g2d31L
Z][O[PdHO&?MEJQ2CWKVDXJP<-0VBK)>C1@5(N(M[V20bCQ,cL<<;?NP)Ld\:N8d
<PJI9C6d;IVC\(:#X.aWJ_I\ZcVNb#@,S,FNJ83W:4dX5Lf+-<-G7W3=gUfOO&8@
bI<YEAV>>GV^P1?bZK&P,S0AQK08C20D@2f^0/KF_XfGM=TK]/E]f7[;S24+DPQQ
5Y0H9X&_LBc:Xd_(LLaU,D#g=B>KLKOCMLMbA:L02^Jd1#5@aMJd).F9]/7L/3:\
.27XGc#I>FV)FEb5Yd9J1C/K5]d,&<(=Y7Ta8OLD&6S=f]_W<3GS\O:/F?&4g/6(
S;/KZ\5;f2HccON#ZdPNU6/2E\Ne#;84:S7Mc3P#/2@VOG)fB9Z24?4W8TQXc^8c
D7F8<?/d@EaQY[J2UePDaYPeV;B,e=6(4gP-G,8=C(GOf)VE:3H@A+OH4g5Z)C;A
+X2_3DgK?E^U]c\ebVRV[0Z_<f>@IN7b>V=]Y9]4<JB52H<b8SO>X_Ma?N3&S#TJ
C(R:\Lf1,X3S51g6DJN@d=VVD7[K:SW+YfWf2R.2]-Wf-9Y,UI-KF9XJZf3X9K(U
[Y=8?-bK3P7#].<?&EXIBR^R^)10;Q8EWXCW[W6Ke_VfVF[;K-S/EY7^I_ZGRGJ+
M>NB67[A6]YEZ6B=OdQJJ.A:fB^5VEM\:G_^^?b?[f.AgE.80-\_[)82b>@.gX,8
eSc(B.ZIU3W5gIPM.12O[M4SYKG?3<Mba[bSa@.=9@>E&M:VA_fE[_:?],3>),=W
OBd/CI6G0A>\QBN>DHX0)DQFO?Z@PWM+YeB#P#HZ@[e/dfD(:SV]3]VQ3#g]<E@+
GU3?YcNHKVEGB),VSY\Ta79a#P#=,8;2Oc1;RU<I<Y\[bdOF5YIbP0_<LN_CAIRe
9Q<-eY.^/?>^;?DOSX)bX8@K:?966#S09]9EC(f[5H_T(@IL0>\a@[=HaF?26KG2
1JbA+]B;&.f/O^ebJ:Q#&SdgEa7YGT3-]UDD<>IgUZY[M;XQJX/gKf9U].,YT)4Z
C8gIN&##&\7[eEZ70;QHeMEgMYX+Ig4cEP[b45c06=Oe,+,&:ELW_NP5C,A4FdUB
7e#2487MO^3.&JYMb?ZNbW]_13X]#&_Y&&>E3@J,f\Y7H@>SQ4?PYdKFWCT16BbX
D>?IT13^Nd@aHIB8d?H=/^L#^#\K=B^+Hc5bfI)LZBP=a2#Va)KG]C=IU_Ebg\\T
FBODO5#4OKVgISZ]I\P0Y,2IVKUc?8?d0=>K.SO8UFE_OE^7-WT(bR6NcH^&1fW+
bFF/OO)fD;agc)#(H8>GG_?]HL6;fceTDWXB0]WH@_61IK7Q@X.UEdVQC4PT\Q.d
aaK/LPAP=)(\-&4Xa5?)X0Y@YIB].SZPQ<bJ02UF4FG(3]BNcE,N;,FR,WK[fZ/)
Y:C0LXKe?D>A2/N_]EEd\7,G[MEgYRWc1Ee+Z[cZRL,D+,2XD4RfHE5\KBP/&6g&
SKK=39#&7e_c]XF,1-,\Ta>@:VH4K+QM424:JGK6Bb9&Y]B^-1,7GEB<4Rf35e]?
)a/L^)7(@b,f]\^B5fO/JBI@L-/0>NWMYGT#X^G+T)=?NFc0Kd9H/OKTD=G3U@7O
M1]TG+6cR26:;J2(Ca2,,84J]=ILTPD.b07\7>>\F=,O-D)ZJ.=W\)(]&3IbdDb9
^-JfD8V+771;^IGX^/-FG][^cE]aJPS9_),_#,YW7K04LWa8OV>W#K8UP\=geGVQ
NgTK^VX^WH:TC\FS&/=#A.;dS(Mb_P<G04L9[cZ6H^;M<_<767aA>;+JU0XfdOIO
8,@D_EdVT=\F44)a&fG@TK_<R+_>Qb1+>3DgP)?4DA8;0\(Ic[9=UC/J._[RbWcC
#/8420],Ece9)>STP:?--#b7]CeU+J.@FVPTdd_gZK3<[)FU(K1>FH0>DX\=8(YA
B[=X<C:c(^/Y9M7VZbg/LUVTAQgN5N<a(&5Yg?bM5FcL6=8=>LH3@b<Q@-ZC5ZeK
RE,?N?8?U-f/P(DE>f?^?L3#U&99NXP<I4[:_^NeWA2E#L]2AC?P:)aKRABG0.X/
g9ZfDD>7\K+\QPC;/E:ZK:6PR1=79g9T0]J1DBaZ@;SL8X\Z2DI/Zf&e,A7RV9C1
QP-Z\.I(b:M<]b?d,fA<&VO\be,@OUH[C^I(2_7/IY;SO+Nb:aVRS^BZ&aRU.eNW
^NW(]F+<gSfKU>8(QHL:=RG(H#?^H6VZ&cD;0;K7\SU#[X8;07d/fYE6DE\Z1c]J
eXD3UNDPQEF,1E?CG]F>#4&F:Tg@(W2:L./3RK/>>I;;FS<M+P)<)OFU=gO&/VY,
TKQPP[]Q\2\9:Y0-JDX(30bbJEP;+9+VF23gM98#HY,1)2S^ROd_U[E+2E:MCMYT
TTa^(#1d13AaCL:@XM7XVM<b)KP\U>ATPP.A<KJK+W&GX/<#N8A#N0_#X=E\/6HL
g;gWW_1TQ]=)A-)bf:OBOa<TK;6:5.a2cJN/1&33(-=:GNe[:,6KaW1AJBUI5C4;
S.C))82Z#MT(b/6F,;b@N2>FRe04=X?/>0I=@#2=fVaZ&b@#=(BK&S4F6]&=O^3)
\9L[d=L-X.TP?.4,P^BaaO;C4e]]4V#:U(9,KJ0KAF=Zc4D_fSF@JPWJFP#5H;/]
S@=/76PEUdgXN:(3B6Q3&CEOc0P@QAIF?_C&N:;ZK7HbH5_A3JOSNA(+<N=T@T#8
;JgfIY=W36\<LV-+.8bORW4&<R8DI(<1IE0JId9/<FCGR3/8PDE<7d_D^^W)+<[R
.Oeb<N2;1\f=<+^=BID/\d0<6Y\Ja=F5O&NBCK0+AV<47>[[Tg90>DWV]&06GJ@2
>6JL?6MM/4#>0K;ZfcANTV(^,<;#4:0JRg]B&?M031(;>CbAED1OcW3(?RS1?9_a
(XWc8+WH1gBSE61>F50_U2A3CPG:B-+EbNYN&.5ECEPH_53T125ARBUMD+@<X-.>
cG46_59=+f0H@=OWW?7^E42/>MA9>_\^LYSc/C@);TK[0/A(6ITR+A1[)d@_HW)^
^@<6UN5&&GQ/C\ZS]Hg;U<\B]:2F;,bf.TdROU\K?I_ORgPVN#cQ.+:+fQKWf(R=
^V>Fa+]aGGX</7g>]35KQGgP:A_4D+:>.U]Z(V&dB(NY_37ZU<6I:/C8VRcbI_aE
+T(TCb42<P)HGYEBF3]_HTMH#/EZHdaMed&U.FS3)U/PY(a>BYJVX+_JN#9UR]Z>
TERaf?X)?LV+O-.\I<#O2QR9SROI01Nf68PW)I:SEM0^W>=ETAY+OJE=Ub-#aVMO
e:#.2e7Ub>JIFc[J9]3#[3MC6?A=A(\A6JP[]7Eb[]Q;K5gF/L;4Y5.CX]TA<.M7
5A1HQ1=;CTD-YaZTAUR=E<&95>AU_/:_/YDMUG.IP=G,-^9A^&7HCY+0aY@R_ZM<
0Jc-L^<.aA\^6?ETQ6f;eN4JS359WKBe7RT+HAQ2dcB5gB<#)d6:R68RN]PKY1)\
H6R+8&cff(cJFMWU]S81RaSQ<CEW>8a@c.S4362^/H5+>Bc3:(Cg=N@C.\]93)3]
;HYU=VcXUHCg_)LX]MUY(_@:Q@@]=L.Y-6eg5a/1SZ<ag0I(44J,Q#]8[:X<9E?#
(;)(72@F[:_2-;gW)c&gPEQLQA1,AKJUf6H@LFXa-P[]H83V2B@6T@P^J-C=38Z^
V\@V530Q3@P#59\>HG4AK2YX7,7L?RH?AJeVc0KDdFOI#9Y#22DXSA#Z</)Hb&G[
K><W_4GA.f7&]aa,23A+a_;)f#&V1?,77&3LCZ@Q[0,^U^d8<L/DU]E)IY73M_eZ
^=F=YNR7RR:9NKBfa;JXQ69[-#2WWG<3b;A<@H8(&#1-N4YJSO^O3:Gce(S(2QZ5
B7WN)0)LQ?#Q.gac]_6_R_-g7=RZ;AgL?P=[#8A),G2.>H2J8@Qf<#?;UR4KC4A(
=\JaGD(IX;)0+09+.=I(86Db0e.@8edAc1YeYOU\8dM<d&R_?KU^&IHU2JQ,/Z?a
IXL3EI^ZU^g(g^Y^[88^=O<G^KI,RD#S>JGb74\,J5#c/KHR:,X@-[7d]fS;)NM>
]?-G/&8aXMZC3BdPeK;aAQ@eD#d\1H1:/=^F<9;8?Z]^O&_Ge+_bH6M9d>0aYdSG
2LcFL+T6gc9,T7AD#:[,/@G6X@0S)5SbQ/#\Bg>WaT_<AO(cdRQ,GQEcJH3]G6<1
@@)8</@eMA9I&X0:E\bCFCEV9g8])=1;TISMQ866O^LJ=f=WNdY?P=NG_g.#E>Rg
W)U+c(N00?MdXMK[d#=NMK93JSdW70=>=#@(#dS2(ZUSQ@D]CAY&10FWd&LJ;41Y
@?+8FDI=UC1,gBGcfWJ\GLIY8Bc@<Q.].Ag?VU->>&ED\eD-V\_R>:58]Vb.f(a-
^X+X0&&f>V>f@.;]O4LcYUM<MU)_K7<4A(e)>E4d7R;3.3JKCFAdLJ:8&#--EQM.
Y8a6/a8ME)6B-WLI:-8VCfQJ^8cT<Q.=ANC@DN9TRd7=JEVF/-=.O;aLc@9X._=b
3N)\-5.UA3Rbee9Gg#I2bL[N0.FY_ZeZ0<J6H+21?7CM(-]2:gH/4c5:C6NDTZ_6
G?eBgKe?dR#>Z3/@dEF+Q,7b_1D[cV@^:GN=PD7<HB8M;0DX:6d1K^&4J2d1K<Y,
J@Y-BXbW309Z@)DS\Cd[3#1S#b>G1^1H<&S=ZTG?f0UE6PagEZ@e6W2BR8B7014W
<FLMDY9^[Bd54gO1\SCK+0=MS&8O<Y__1,Wd+cGW>1174LS-XB[_Dg=0GGg>@FR4
-((&H?Ab?AELM(VQ5Ze>gVK\(N+OQPH,AR?+Wf9Rg3]Q>GS8ZL>e<fDe[AY1SZ8[
aLc).Y+b3P.)246:H;Q0+cQY+_7YIUBE2GHacf7=;+TP/Lg^3Z?8DXX-f93@76&]
HdFgH+#.=La\S,7bgA\1;=g_8;6O^9+R4cW,3LS<K0PU8Dg7(&QC=-2.R@-bR21E
[1H4;@Z]6\VLFPS,gg^U3]>eUA.RO[TB--V\I]_)B0c0<::\dJX&1H144YM9I7K<
[#19JZN:P+C82F3fY=:4V6_a^JD<XFbBc[T0V-58FS/_2YQRQADBcd:^\<:A423<
[^Y1C8O8/E^[#743Z<RM+19L)Y^YN==5;d?1[0O4N7f@@LEQ[>gA0\;I9Q77cP-B
\JH(FO8aH/3c0SD]7H13[=C^9>RL#_D<?12JK5E-X(MA(YED7C51)T-fC+Z8fN^6
WC]aaL83CGaLQ)ca6I@N6a0\8)VAF(:@&[4aK]NgNCS8F:XB+--QR>:PW3=EVODe
G7>89+f35S[J778=L],CB:]:1SUS2L/PTKfO-EG[G56_=d&<\Z+7<<&>-R\GO#,Q
8AO?0_XOP7LPcUD];;GZT^1e\L9U<_,>[@.EH@42=0L+;NQE>\]V8=#J6efg9F)V
gCX@.>Pa9ZG-T/aO)7G2FB+6N\>;1]OV_I:.LW[KKHEd.@0eS91f7-4MR3L^(Dg5
PP7fR>UUYb/X#BQ8VO7[FQWI0]O[bfX;<7[+INX#]=gV@M66KABeWg&:&90c_fM1
2aEcX5OECRD]_+G5SKZ(>+4Xb+b+3[S[UM;LbJY4/DR;VKQ--^T+^XS^Tc.,5W.]
PT;;S-\g^U<g?^.TBe3a7PG/^1^.b8gW8+#HB2LBVNHf)PeOfU4@&TI3Z=8)J[2U
>QgER?8[BNJ=VJH(Ga#E#,JP0C8>=+@W7Q9FY^X8g27AeI-0-[T)+a:FLc/+(VcW
db+8O-G;<B..cW?)f#UP1dAYZM>_QZC6Ac64K(ZDf<_<E29/I>ee29b@+;5)bJ[D
_:LI1^cLE(<=-eGaA^SFRVUc]C0LP8=P3/LBX/BaLAdU\CbP[T32^Q:XbG\DI4]S
UF7Q[IFgA-5=SA\)UKIC)FSH[;5Xe7+[I[4Q[_(^GbfW5U&.7WW&_OL988aJ^RKI
G#8B7_R74_1UJT/_KfQQ@f(]8B_6,_]ebgYaTe#[<&<.PY.:D4V3+8R:T,#eMag8
72aAd/OfJW(-520@=^D#BY#YP1J([[5[PUNP+b/1\H.U#V75?RMM\NJ[G+@W](LU
bNRTTR)IIfdWbJ]O@@F+e4aWCeP.U[61)dI>L]P,6fBM1(ReO9Q,\>f&,)\Y;[@T
4H/4PeVT\)0CC4W6F\C=JO5TG6)f#4^#KS\?:UT9)cVc5:I70;0aK_C2d4I6G;ME
Z<Qa1a6AeRMF:VPIJ0/>5?B]804?6g8EaAPU;9H&(:0gB5c2Z6-[F74@G@WVKDU(
1ASO@O>708\a3EQ]3K2b_X-XS55YYR;YFH.=7UVN3_GPAVNPRJ\0+CBO30YR&GeG
f4A]ZaZ<I(R.GP/8;#V)f32,R;7>Pf4[^]8@@d1<N_X,J,5g+.c\:[cd.>;.TUPZ
_d0^@?OX0X4Y@gM^7U<S-Z17DC<XB,_dT\SKN,4=a>^R0/P+X;::@=dMPH26XZCS
BebN8R39,45^RL+66&Ac<&O=#?=RM2&HO/LLRR[K=B6+SZH268PbF+TbALSNfE2G
PX;9G)X5dOOOCI3IF=^af/@X?Zg\/1X6.7f&0W[Df<ERH)QDE/OTG?g-_<X>]0eC
[@Y)>/W57CON&\Y3bKbQT]fZ?(Z:[BL;XEV1RT\WEPD;><#.<XEJH^HQR9TbBT&<
Z88@QE5&TT5>#CZ0^.a;(1D3I89?IVB+S(UaJQVQR?<PC\_EA>AM&D6bK#08,V;8
S;93Q::_a](dL^)ac(aN.)N78(N<C@74XLU@-A@EdfPU1/GV6.:1UHGSU)ZTV,B5
Ga^a>^F4W8>gH9]56?I>e5X39RM4AA:@080b81e7b[^>KMYO_7,I0aT#KZEAY;D2
93D.gST57[IOUQ_<R7@\5(f>MQA.N:e_aS+(9D0DPg=T88N9P/]eRdIM>Kg?1Z6T
P//[TPCCgW4V9P-SbH^7OI)Q1-;HQ+5D-D&Q5D=<TTU@2KN_@[&9W,SVW^B2?)#-
\4AZA4LB0TL(-ccMQ/_2K6OGX7;FKO?>@/F\aF-3aL;5bJP?-Q66N5EdU7_TfX=I
SHd(+I3/>;]#<;CBBg+UN1<ZfZW=+[0RX7R]T^X_g=e63Wdc1PD9OA.;X?[d10=O
TQ08F?-,ISXc9<LAFE#DOX>b>,VU7-SZPdODa0-2@Id8F@@Z<JJ-Z:X;XOIGLC1c
6[ALK)9)SH/1K65d5F8HPGeE]/8NAYH&,#;,56:4;N12DAYI/J70RY.c-GAcaBf=
2;/S3g4+Z#+HFM/]1eaU?3UWH5M&</EHGT]2/3GbZO+J76X-8eW_C[V=Y>2Qc38)
YW((_))U@TIg(\;1DRgIDe\5B7Na:Ua2A=.FF_KGGR-WNag20BGY9G_<fWWYeXWY
<?dGEfVR.S;f3PIPZ(852DFb>^ag8Wf-(FU5#XDf]-D[_J1IA_3c,ZV+f:1K[KAd
T<[#7\^.Q]0^^(/\NE+>8F;>VRTaMZb4e>,ZA_A1;B,WS=Ge@)SNJV\AI_CZD4N>
UIgA0aWAXb)Z:8,^ecdVg#ZBFY-cf4[O0C:(F.VaC9HXI>NFH2b09:Q?^0ACE)]M
N9&ZO@Q&C3S\fcX/eC9-gaL,e:QQUQ5dYVBZ3/Xag;e4\=VM+9A;YRgc0#60I9.C
(90DaHU&cGXCaPJ_O)-.gbA,NOKb6(EfWc:_(bP<D#1_2bE3;1W^Q#D:X<):cFG^
Q5K3bLg^+I18VEeW9dXL-_L<>9T6Ue948J2>U.]O\H4T]8VMQB)G@Q3)Y-9E64d@
+)1RDbadP/R[-4g-;+J.RI[3>I&OFGEPXg6.Q[<G[(U>T35<adFM5^^DB^?-AEKQ
19e,^29+fd1UE_FVXC@Y<a4bL4W2c?RMN2[=DefY9T]BO=N\bTP4YD][N9E(#=)Z
b/?=VUZY#YOJ58^VggG=J47ZOcMA,bCe5<4PU5+gH=:Qe7QNX<+K,&,CD2Bg3BOJ
F=)V@@EURR?-^G2-G-TTIX?^d[@7>dS+Wa60.DYCUF=0S<<2YD<(3b,[--a85Ecc
f#PP_(?.TBOgcF&YO3O^TK_BYT85Bc?NW^^+gWX)cC62:1(X]OTC+-:)5<P897Q(
EB=;(GH)Xb1@I[RA@_e:<Oc)))#O\9LD4F>f?Ff(MPV7.7I)7)==?\c[0R2S.X,M
[dE67,>?f2_0C404HLc(=KO+VE6d_Q,@4D:bge)2e\P2?aWNBB((ESPg6E4Ie#P5
=9^7Y];]9SNV@[,M]He_LTLWXVT^VEBM;baHEDQEb2&1#S<+OK+,7\1Q)<d\1LA,
6eNT-.AQOV\eQ93=a1OO1_=<Pb@d78>V)_KTGS7TEB1.?QZgY_3Ye2Nf_F=eVW7Y
\6W)&-G:UN3dY.V.Pb)F7_E9CS3T;IE_L)X)_A&,e0\Ue/b,DMO>QDA2J@OUdbaK
[V&O0&d.4.=)Pg/ZA7d9_BPUR#B6(XWHWU8;BN_DKe/C)[VPZdN[I>5L<<XOO^()
FH.;\.G0TBB4?K6>EC>G,6=&AS[ca6T(c-S+E62WNY@BSKJOBI7F-5\-/+&N-Kf+
<+gNX7C6Zg8.eA-ATWXAc6/H;)YB@^E\_G697KbSdCKd]6a3MXK(R:1#3;SNG&\=
LEJ@T<bb4bN<R\BaBVDM;_AF4:#D:bSC<BWBME5+\)LN\B<D682Lg:e;N+J5bKH&
fPB/VQ(=d1CU3f@/-YF4I(6e[Qd_J?b=;6L6O@MJLTOQT3956GTRUa@U_Q.&&Lg\
M&4bY(,MeWI0(Z9I&)W-V(.=I89=fW_9.9W#Z8<[]UEYOEO4F/(\.?^V=aOUM+K;
b:V@3Q5cE=KN>GdNF)Kg(.680H0/^(+SXW]_X9QgURe>EE//eG=9G,DR7JHTU7J@
dF-<#:URb>/T)cI.TLL@c]b5@J,6FIGgOV[JbP?:9:Z\M27#ZY:e?L;=N??YTI1F
Gdbd1[2R6MQ8?6cc-Kb6>B><e&@2KD7IRf2feM07FFMXPPMe/@VCcV[1dKCO_YB@
.<P>N,&Z^c8fEY#\g\.)RDI[W?T0>3c1=F8g&c_++78SUR+Tc#VR<M<3Q>N(?ZG)
Se&4K^_ARKJ@/HM:]UJ-VbA)^J:VW)/+?@0P8)5)\P)YZfH[M1@K3PZZ&fKBa746
H+;_T@fN(6^UCMZSQZQ.80#aI#bF>Rcfg&ZZFcBX71>GFYIO:PX(F7+#ZR8Q3/W#
e]GaPT1F#H4XgN[E1F_4gb@BT@<KMB3#M9Q3Vf=LIUN&=gd&_gXUJ\NSR>>C_;:-
f<72A,Y#U_NL0G/QLA3SVf,]GD+XUK49aUa^9#PP]4P5]Q^ARB2b0B(.I.EH3OM/
3ZfOH]Y40Qc9#Ce(_G0?P0/NP?6cS+7?aSV4JD6bcJRX7WH0EU>@;cW#:(?dR6aD
TPOcPXcVPTcU8[BM2ZIG#LE<&HXT11/&U8P(&W4gRS&GZ;=ZfP&(;8,,0M0b/K;V
:/)UV>QMQR3R;Y3N.8eMS[gY?VWI?J-PTRMbF<:1PTO9)Hd8+g(.)9)\F2b]T2aE
[c797_3,)+^UJ_?d8\EPcdA2[-JDAJ,KeJ/N6VA8#OW9408<ADSHZ:=:/Y)C-3HY
PU[3e)44HHdgFR@gH2Hf-g3@^2=0,S/ab=1KJGG,Q8@/[+W)O3#\_.B1Q59.bE=M
@WEHdeUM(H3,/c<:B8L.]V]0R_K/Mc6#^S6/Cb@e@-TUQF323VP983g+COPZ>K4c
Z0c7<KY3R@6C,N/OR5]#0]ZZ8M?]e@a3C(_UD(S-9LOgVa_ZaP\g>1Z:Ua>K#AIe
d,56ZGNJQ5ObBQU9BA@HC>6LEEbSKV,;?F4#MPWSVSgg0a(U3@DF&1YIDQg(gUg6
-6/)J5F/)P:OY.QPHX+8>L,/>IT=GJ@&A<1GCDCM6e8#<3@&AI85KR8-30C8G:Oc
a,3KXZcFfB(YaZ[cUM=)/-#-./Y3CH4LPS#8<G>PC:=4^<[[4R:89T^EL2YH,&_1
fDLLC]3RE8,;FJV3[>QT9?2-O];I4T9-=DL2b_NA)aR@Mb508BF9M0\67T[+4>0Z
),R,2e>5JLVS@7_<]AKMKNgVO2(?2]@DCS;P=\,#cP2I51V[Ee2^YY;JRWe>,QG]
L\@U^e[5AbfR:LV?adENQ7YLD,>0?;FULf=2N)d+/J&(_g2aeFeSKFg2P0N0.N4d
+>+)?5J<CfR]W@K3dbD<][LT<8AQQ@g]Y8U(J5H_U6M^UaR)d?1-+_:5=?3GYQE-
6^I2N6bJebZLWJ,N[8Ka(,+LW,>:SP))c/F<4QV9;71/?F0;,D6[cE:CX-bE;51_
CV_1+-G[-D@3>JFWV:#,M--7Z1VKOD7?WQ8F:+X++>+ff2e++PT(3#bOb8LV0(\D
Uf-=IK#.V&E^:P]I#b,-BGCC^P0ICD_Ge)5c,fA;M5>G23fDNUU9/C3;\)Bd+7M/
3M,.=MIQ^7Y_XB(1LKa2#NNNZ/8g-gc9)(97?f>YaL_bB0N3dC:?:?dVU@:X@:SM
78FaQLN_dWHSR579O9I+(8\BZC74XTE.aJVNS-6geZ11@30G/c29g#OK)2EKYf\C
B4,^95+0B2.@@3@a93eI22&9>fc4Z-=Ee]:=3M,7:#3RG6GgW.)?2;56gcLIQADJ
IZR+(O&WCW8Td)aBR0Q/-9:ag)H?<-R2FP9S@W8K>I0cHgHV1WN-3d<FPX0YGOW^
1a\aGY).ORU,\91\00-ZGAGF>6)(0PA^=eINJbQQf11-PMR<R,D4dD=CJ^PKOec,
[#FNba+FPI94?=d>+7]7MHIRZB<I#]94E5f[RET5I7_B4FD3PF<HLR^T2QI;3;\:
+Oe;gL5GI;Z&Q]GQI9dW\26S+OGXQIC[(#18E59YMO23X_6@fM@90L;9X=e4b;)&
S_T]/T/AY>():CA8bG4_-XF)ZRf]+_De<W5R(O6O<O9bPAfgP8/5;9H19)F=c:1Y
D<R)g&b.EK_d6QdRA@aUT[cG@0BI9&)\e-(\P0U3SQ\dB0PIf&5[4Yg)2,fUA-O_
9V3;C.+V[>5Z0)-(EU/#OPQ1T,cSBIK2CA&cN(GJ.[0;EB#YJNF/=>9?KVHaUNfS
7R>f2GEMEH+8/3E-^L78@[eF5:9EG,/L8OK5(/\6L@IGGYUTTNd;(8=<YZ82JH@)
([D?H&QbA8V3^b8(.BC8Q2B,7\)]:DMD5HEID4I^4,>::6)bO5N+K]Gd7-Be8&,=
FGW1I7)Fc?Y2e\O,=7Q_H_=S,[\<bfKQ^4df]PA\5ORDG;O^MEUH;RQ3Z8E=52:A
L:fC/Z7gM#_a>LKbBg2[R_8:+6POUY:6QEKG[<;W<QE4a12W?X>f;P7<],EPKaS:
HQ=]f:@FC-P]Q>AHP3[Ubg;;e9MX#5.caZ35<Y?@U^dBRL]=YHWV5OP9g/8a<7c,
_eG<_(K63B[Z7,T8(K5:17RXS\Qd=3d8K=c8BP--FDW-b,F(K#3c_VF:g&OFC=Lg
@&c,=RH&Y.VN,V.7_(6&7QZDefF3)B]W?D?&@E7<#49fF_2I;W=/=YLbKJ]O4?93
8aZZHOQ=\gTA9ab1,WH@C[Q\6TEIUOKZ5gOc5DU;(3]>bKANU[SXC@K[g2#F;7.U
TR?JLDa-bW#fD:D35KL97B);.,)\@?4)P#/cHd<W)^H1W_3;D&XA<Z2QVb#De3B#
.>+@J@L&4YdZ10[]=AX9[dD&A_S?9UB2..52+XRN\,1S&.0T+TT)X#7_&QDR<^#9
:gC[):5G27P^^,Q6A@;RIO8gR7_-e#GdEWLT,Q=;1,]RDVJYL>9F@#<4YW7:=++c
DEO1a=8=)[c/]&BH8_a#20^T2G:4D>=1O426#P5IGeaE^fb#-/Eg:eRf6E/Q26R;
7f_,HRIV2<ZTT3+6M@,9XNA7aB[^([<6(Z\JN>I=URfB(JY#@;-MF>^K5W3):E[:
QU+P1\_0^8@7A,<3)CO7?Mg5;^@<X@Q1WfVQa5Eg+:6Z<JcJEPcG(]fe>+BI<ab\
[.D05c=(8U8_,1bE]AP^[+H0QSQ8Y&>cfA2_UU(b.:IL-bYUVaTL.C=A\PD0P)f9
>VM_]K(:7QAIVZ-SMgWJg<PY#TeX:8QU72,>aL14-fW54\ObGe<P_J)J[-b2HVXJ
WS]M<G&4B3Z>(D3IC@DDN>?WV.1cIdRP)>[8MPGC5LZF6)?XL\.6K0X#DdXQX[bD
=WaR7X-fIWaYe5UM^0>-8IUeO)b>Oe+:RHPIP@Q>Z>cd5S?+/T3E3^N4?[7CeVH1
XY.EMHMdd]]#V1I.924H4[H<=7TIe]1b@<E1)LX+BV#a23^&F=YN65<YVLS7Gfdd
f]9M@g(I3?I.?BOSJ]bZA3HYJ<W:]U=ZHB6R5SY,f:7#_YG4J=KIg2HY0^(>E9ZM
WJX/aTT)ge]WJ7)X>aYa8_YZd6b2+7R>,1XZ#6255PZ5=bSWTA@bf57.-[#_g4\4
O:^&,J=g30RYT9gf0b(5<\O4L3NF)SQLBJM\@bZ&bf_\1DB.^[U)T=IK6>L/[?BF
5g&_0;-[-^AVN#ec5[;1J1c;dZ?C+HFS^Y]IXYbU=QP.gG62RJJL:EWUWM<d>J6/
C^NTV=JP]B8E_,-E]DLV#0HLC@W[G>>YY2=C]KbQ.KC_cQ:G=8#SaF9g@_+?LgUK
(9<@U.+D3T[7@A<e21M]Ge@eB[BQ\+=9fS_L5D_#aQ)?59,WE]XFKA1Z;-MB:;Cb
ZOJ2PE2\T+B./I;6_0&#<>^VS]CBWJN[P+=b;6.e.F=^39=G_;-H+g]B@KJTd3P+
(QO7?.(M9-/H-VdZFeeSVX1>V/PHW_),@=0=a2fR;&OXCJTLeJN)Bd^4><a@fOaZ
E+IA7Z2Ue#O/5^DgTF9OQNb)ILc)F[NcC-U^7R]:7M0]1?\3aB,IVNc9)CN6f7N9
:ZPTR?g9KAdc>IP&[QdO^HIe6bAaU&5YT_VWCU_cB4(46QBS1A1DZJ45CCDD[144
edFaWOUI.RU:SX3:=^E,Hc6:W<P1Tba;U:>?<M3H)3,F(;a/PBI-;V.JN_+cS/1e
DHB+&1G-/3L)KI36)E_WVa(3CgSJ+g(ORX/>Ma1BcHc1Z0&S4:c+]ZdOA\=T59a]
N?Ee[=[E91UIU0]TTV&M+gIaaa&,.OEdO>.+NgO0/8cbdaN1G\e7P>&I[@XTVO0W
XB:A#L0_F>b,P>gQQ_://&LVYFNgZ7g#E1De(3&RcVC)HJbQAFYc;4RU5H9/)WP8
9PX/[M27?dR3?E34f]L+=&UI?_\Y<1P.BQ&9f-O,7[,^8SIQ;@06PAPD@RE#X=)=
Z.Jg63aC>AOd0TG351E_N[?;+GHce)464MN7fcfC,OEY^[.Ad\:QPbQJ8)P::7K@
gDYSOYTSTS@1M,NDB#D5>1=&^/H2J;OQ1;>Z<S5NU.UF59Z_TM7N_>HM-eUXS;Ia
RZa.\\W(\HC34[?[+IBN<8<N?LVaL:.H+_DEOTDB.BZ:&8XDebHP>-LB=G_gVe2G
M-.XG44(G>,+>KLOE[XHFX>4McNU4F)M#d7=^LA7?<EK8M_1^[dP_H93?55,8O7d
#.I5JXaW.XTK<]?B,;e-c[c0,(5W=JHTGD75>KB+-9:0&5NHC9[M^0U57P^44(/d
L+<_=f#5<8B11gRTK;6OH0L\9,B7D]eNG0_Z4JF>HCLOcB5VcL&U9<7\e2c[CPK-
?3deU:K^]+)C/EI\ZAPOQ=(.?>:4<+_1Tg+e>CB^8(]#CRf=7>-XELBN(R?1=E#X
?WO.-F,2>WB50YC44L:T(K^]7E2HDLaLeU,=5HJ.9H[6Y:ED1C\K.WgDgL&Q1UX&
&_G:##T.^9g)@=,<]9&gZ_d-#+f9cc@fA-/[.e;;;0#S=7GG2gSX^W9-E^9S\@CI
d=K@BS]#\aG63eaHW352T/PYDMeg:-9;\YORSa5H>K=1VbS7Zf]e\<C@)BSY9)&g
^EZVYEA1c@[L3]F8<:MNM)7abU+6fVAEG:Y9WLSZ9>ZP7IeP&^6eRaT(#5c\b;7e
PFKb,g-T@4=K@[&B986fX(<.D0D\X0BDH2?^R3@XNXIFM6;9b6B<c-c;L7eQ<<Nb
2O,U3_gW01K4]1Pa85gJFQc^D<8@Ag<UMgR+HDg=H7B6X_b\XN?JXUCUg#4Y0AdG
YcU.W+)ZD:9a[1HaI?F(f.,XJJdd<7H<d>C\JC<=L>;gCFCIJPC-1AY\e)3&7M[c
:?ICC>7;(L.VS(V@,9=.D2]H<;=U3+a)7/]Ie3C0X[1P;4aKM5SWH2&EZ,8+10Be
;_YMeY4Ug.+,4W?e:Ma>:f3dW&#S^S1dI4QJWE1:CVK<e3V3I5gHURcX.4^WN+b0
2B6dT2IV2WG;IR>;K<-Y6<K<IP2bY^<#f(G(Ae15N&9bTW@);eD[Mf+Ife2TB7CP
CWb0;9MJe))>;4B)KUJ.F4HNaO+FKFYK6T[a_75aT16.Sb<dVSADaIJaXK2&B-6@
[c)f[ALBZ3XfP4L7(^e[Y==#HJ^9WU^]@ZTK@7640b1UN+PBE_^O?QBWY15a@DK>
&1f73W[BZVV-/[QL4A2Ze-7=+7UR79BB-PV4IVdE)cQ][8,C?6V>/dG^9K9-Z^c8
gccU=dYW_));,,J#K2#-]6bW1(1[[LO79VL>Xe/(;M:=0)AGBRFI-(U5.f)A),7C
R-0VOAUKg4M<\LS?8UA=)?Vf54RPc_7O=()D_6D(e.(g_R:PYU?NMce;=JA&_Ob^
W+=T^.C?H^E49[2c0R]#G@cM[V\N/Ia\]I#XfH\bN?OB-N@^JKT\(-C-24Mc1a+L
6Deaa6PPf-[Q_9WLe_LV,bH[+bI.4PA&ZV#9]U^V5H76e#9H(2<:D<@2A+>/_C=L
K?1AS7McO58ICDIEOa)<16BHc:Z36#e/=8^X]C^PcSGV9#[W+KSU&\:[Fb\:F;1)
KVF[J?dNJ-&f9U?E.>[GDR1_>-Wc>>-W74?F7SW->E@R4RB:72D-SHIH2FJ0+1_L
#L(+YYF,_4.@[B1>0:MHL)65e(;@D4N1=B/&0+XP@KX?2^eC02LL-49,^NAA.G74
S]Dd-JI@Xd)3GbC6b^b/[>;DeNN1:0IGg.JT<,[PD<Vb4ZbZ8Z#Z;JScO/QR-I>b
Z+I\.HRS61;L<H?#APT6-2+D:SD5\B&>ENW.70&2#:)+62bc1S)LI8f\;8=;\W]Z
M=2W+9MK\.OV]E@#b9;6H5d&cSBH?+NNZ2OVc[3]DCCZac\7=,9dCY9(gFO0ac\7
(T)O76C)S:c(9/bO_,^fXD?P=Gf>g-WHV6)4^5]=F2:WNb8f08;BN#2aT[;BfGTg
?G3G.Q&ag=P8ZSP;S=]7^YH:][I(-aH]FSRF1_--Q4g\Y>Gab-MR\,IN(SRQ.44[
g3Q<1]7-[@65M\aePY574c[(MY2OC,7/b2WJ/CQe,,,(4MZN03cAR]B,aLROdKTL
2EJLNX1LD6@Jg)W.g_7A_[&YZ0^K27\NNQD-0&cc,6\<G[[GOZ9DZU+OJV(_J,30
9ICYZJYWSX+W]0(\.&5e?-:,.RI[30eG-aTI=4(,cU^7819ZZT3E;E?X\c(KEXK>
DW3C;0gCeF+7/46(7H]L0dUEG4D.4<4+A]8FH(C29BV49:8_dTLS25&e/3FRb0d5
SEbB1b#<d&-BB&4_,]O?c.CJ53He[6TT]41VUN41B>=a>gAO2FG6Sg]X]QU@GMV(
B:7T_gGE08+g,A^S<POZ7f,D?<O:-,H;,W<#bTgd8b+FR):Z8=NdGOR(R(:Cbd[b
?H1+]:(?Q-Ld\+1UVM,0WFDJL?S#X9E,47RY?#1XH@L\[:71<.U0SSU:0OJ4J.:\
<G)T_\;ZB[G>d_))+9@^U6QL)ER1Q/H&G>S_2cC0U<U)YP9<IcY?1QGW2?Pf,UF0
^[JT5TY[8W3ZPOXK[:6>CS--_S,S8Y1L7</+WZ2;QTD@999FN(2G0D8]_8\g6&Wf
7JAPQ<cc<N46=7@]9?N7S5:I(_:Zc(]6&1d4K805(\EZFTUc;J59:@2M)Be+S[C5
U7=7Q[/PZV1S[cKg?Q2Xe(.f]+WLN[C3(b(OcQAc<GTN2U?S9Zg<]7)7SYQF^.L]
/FM?.83COf(acdEdXeS8CO+b[&8/?::DW17IAAaCeYU0.aGE4?KRLW?0E2WUe22,
Q,W/QNcMb5^?E.9PQ@2-EFE#UI2(5L._)>F=HdHM(ACRC@eO-5X1V9Y@gZSf[TGJ
-U7@;fXW2b@_dF,<2NeI=OUV_)fX9\YQeT&]KS#@M[R5_9-&-_dWVT2S7YFI-TGR
\d_=?RZH&cYZBALc3gD,[S+X@7d6X_)F?Pb?=7ORK3050))e;+EN=0(>OGAe/ATQ
Q)(J;f&TU2b,P4KcQLXC:<(P04cH.?N,2NU(K^#F^\b2QM)?f03+-Z67QOJ3DU40
R^<MC9bcL30O5J2c_1J-L^_Y?0YAP<BZ9VU[4P4SX;3:EIL25gZ,S-JI\P3<RC:a
Q#e\_;#S_L,O>Y4@O[0fBMUGD;FY76P>2MO4V.adJLTEI1M=8A5<EDEUgX6691P&
X9?[<@,PY]=?-?5[31,b[19#X/)#bV=bdY6^W8dERQ?:=ZQ2,F#7(\@VP0U/@_(P
DF?(FVFZ/K)/V-4M.\339cGN+U2<L9N8g<;9JE@BN;_g6W,F2A85E(eFVG;#PBDU
VMabA;cC=<BI;QQ3QKOSd6+7gZ>)1bS3gE;G:KB80.eL//,b#6Ud9G9f299Bg55N
M<1U9d?7(ZSNB(bY#9IVU??81/\7+AE6D7C[LCIcBZ=E9;_UB)06PB=VQ6?;:6^c
(gO8]I?Y5USE?^Yg=O6)Yf.KBGfgY2C)NeD^(.bAJ3P[@5GJ#(.,?2MU\#bb4J:V
ddS]].17RbIWUg76Z^1d\V5NHX/RAB4PL6e;4O\H+^X42UCFSXeWgBUY\a2a;=OT
M7KH[>L72bE8N;.D:a-e\MHEFEL/aa29IegZ]Q[)BbLg=-\.+ARVFFC>\R;9D<=R
OJd+^_Id?U_QG8,7^Xg7ea:,7V2BB&5(MTI_X<TVDC<XYNQV_Da,#>Y-/Y7]3.D+
FI:)@9d(8ccc=Y;(W93?Ma=/R#32Ff\4#-Md]K5\(#5Td=52W+L@9YXdaba.Td03
Q]\,L6195,RU)R6HGE0EU7cfbYcfbH87]?7/,gZ9f?G)dMfJ3a9ZI-Fg[X\M+.CS
gK.Y)@0?LK<;L_dZ\\+39OHAA7YE_/XYFbW>QP@BfFISAe[1V(/e6M/AJbdgS9@R
-M.Ce)V^C_H0-U0_f=0Y6&(aRMQ_@MV@W@M#CYZW;D71g?<655JL68CWC;A+UX)f
HYA3R;,&@&eC4L&02[dGJ+TC_BgFVY;VAR?4;DG3/^GEZD#WQ:K,E4V3DP+8)GUJ
39SfT9JYZ0G?8)?TY8a8<O=>[4/40WH[C,MO:Y[Y8_MPFCXI48T36H>42OHCV3KS
YSP]#B5)MM3gd?^gfS7XX=\@[(GC;8aDaW]B^10RVTfE+<82&P/@1[Z[BU99<NG\
aR.03gR^CL]0QGLP[6=-2_:ZHeB:T:D=+C@<(OC+2)6\1J<c[TC9F^P9g0aSTMG,
B4AP,?//4O+W]Z=9]dcU:U5^^fISOAT93f4g4PV([BIe#gR3=:6\8-C9_)/1NZ^;
BB3M\X<fDRO;&F:D5-4-E:H/57<7I?]/-A,890d#6V)4<;dbTYa_>:cgg_AR.3-D
^V6EID5eB:7>[;LYa7[M@4M6\gO;d&a;-AADa3HOd-ONF=NI#_ZVVQU04G<;(J)>
1CJQ_fEg3Z;_?\^F+X>g^W;(J[N-L./P)?YKTI:MgK:]I2:MJ]_?e@LccRE+I3-:
X2WTV20F^<VK[M36[1OL_L7gLRHW[&=6X@)K8JR.CN>>Dd@^VGY_2.\LWVa>>1EI
P/-g>GaH.)Ia=2.gY(CU.BPC^PfOCGREQ)+26C+C^/13MT>>G5GD#2dKAF^U+MDU
/O]]W&gSVNOUF]J@a605/95E<b,]@b<W.)>5&W1bGN?J3e8eFE5=PU?GQ0ecI91g
9RQT;)LdFVaK6QDe<_I]&eA.a;IS5R&0/S08C=)5@TW((D_HC-2L8L;@:>UM=KdW
AG:OE5c8&a[F//SeR5D:M4a34EP_FNY]<G[C(E@6N\Qb\Y.<ec@)1Tda82YcEK?<
@?KS-K#F6P.XebaWe1eNf5JF;G8a8PX]R+/S1P;./\D;W-&gTUZ=dc-(\S7D-EHA
D341V(1f,M<OdFed3=V]#1e#U&./+44L-8I7BNJL:CT]6Q234-IJG23]L^J@^P0.
C&_F?SZ^bL;/,-U#TXNCE:9HY(LgB7=E)X[>EIE>L[a-68\68+=&B0I24#O_R2/A
EAU:O9?A@TQI^X(IVC7O04BPbS@V&9LbcI]2Sf6F@;&1[D(_2MC<0GKNTa^Nf&SX
0O6X62a90^&YQ1ZD5R^FJdI+[bdOEGJM/aeXEI3)8E#Zb-\3YOHa>)I@XF3I6X0&
><b)_\Zg#VL\g-(PcJ>Y-M+Z]F>gII@g\81SEf&,8RJ^<4Obd03a.b&UgOK^I-@N
ZF#)-4=::_W6GWED=3Q4&R[[SID4fcb1J&F7)]gZ4EC[/2&QZE]E5P,VD8<b)BG6
37?M.[V]Xa,FA#,]GL1/BaI_RcU_^,1<81Vc,6Z@0d22298f&D_gZTI2cX)7^<aM
38(I@5GI,dP7V#b/J<9Q(SC(F,QB4>PPZAD^(F3d,_O;30LcB+Rd;^D,d(dLCGZ/
:28]O4+>QR)QKPd[]+D,(6-.UeK6b@e49HgF(d9S>+eW@HN-NJXe<F.CPd]6g44U
9/EXNZ)3YK^XV-OSPB&>WHQWCEH9&J,W+/=_gaAAS)YPfbV;&d.e\QafT8/3KB,C
XCT<?MW7.3NY]AO.d49L#2WcK_V2E0(S_F<5><74(],SdT7c@6]g\IS+eO?_(IcP
^B/JM\X<XQ7S39ADb\-PG8g_0U=#a9Xf_<:9f=S?02TQDB/Tg@O;/cgZ_G>HMEc?
#b=:(@NHH_,Ze04-+10=\B1DbBFJIBJZaY&3Zd5JJ4Pe/1HWUHF6F5ALdHY6):3f
FV)fC#aREe_>G7>Pe42QYGFKg=]8<W7AXQ?gQe]K4f9),T@^-2/&42#652]_]6<-
@eEV:IDTNDQ_J.7??/-/De_4.SXVB^D?SWYVRUK+B;Mb>SW^Z_Cf-_Mca0=^GfSA
\B3[=fB//;15a+0D0VR//Tg1EH]9H-?8TFX9+B/9B7V^>25A.PObA5+).@A?#8aC
aVEEXNM-)QI]OeAZL\Hb#&?4[4<5E0JZ7;)#61Lg0AKD1-We_?Y-+?KY]KKQ3a^^
/#8.RKI3dRE3Y=^g[[^_B)NLd=ND4V7)5T,3@.KG8Ie[F@KA.F44bg(E4M_PF;1;
VHbP;BC[Q8\^3VLZb);cSDJ>CA(cKZ>4_85G:A^SI5S>CF=)1K(/_:#)K+cOZS,P
47<2:cNI.2bUgNAJ(,&g9]R1;Wg)Y?&-[/4f3J5LG\C,g7.;\@_#/PF3YB5INE1G
P_HIQ?B6IJJdUac;]aI4YA<F^4@;4#&EYb</H+W5&0]/#M&/>84Q<[OV6.+(TP^:
T73)#?D-\)dS)WdD@B2TVGV\.WAWQB>1S.6Md);9IS1G0fTFU2eWUZE[W#=LITgf
I6\XF6?,@L7Y[R=(3..;.Dc<CF<G;2cO:B2QIZbZcJ]@GE?PRMGBWJ?eL]./UbaG
a[-AY4Y)UGLI,_Z>>X=NO:J=22F0(KQ37#VU2:a=BYFYN;H<VC?H5,JHNJG\(02?
_=c@BbF;#=SHQJgZ_dQEP\=J,d+MR/+AJ_4DVaaB173KH0=5-e#gf1<4?e_PC):^
N\ca4O[AU2<\eQd[11Vd-V?WZMS.YO?M&OX\f:)Jd:R]P\#LdDZ/[eJQ>?9BgcDA
e(H@KJ++>V,,^a[.Y3+WQC+5BJ0G2XaF)-BHSf5dRX<bb8/OA98O^PG;.0-a1O[.
0\IL?cEKdAAQ<I7GT082)X6B1LB0CebageE>/9/[AQ;GVAMRUc4c3UXgLS+(Q+c(
&-HB,7=7)dEg+\(_6HE=X+O_c#eHJ+@UQa0Pf:KX_I?U0K3=aV@^\L=U5_:=9BRE
-PBN^NH89MU4gP2Y)b?Z+T?EAe3@@99Yc(MgG(0,S4I)DZ>g+\X])[gG>@f/J(g1
+VE5>\N</HE11.dO2]\=J8APEGJcY@J/01g1/9\C?Hdb]L.e388Vb#S=N--KQ&L0
PX;P_O+2e[/T?0C?LL6H^&OZD,V_>,YUN7/aY+9;T2R0M]@[/bU.0>[bbg1:==>:
E4\JI_(U\U>X]O6cUaFQ3ON?J68+A(0\2JC?Q2,^+ZK1a-9Z)bd\1#W_g;H#RL7@
b[A,Tga1XOg)ZB=8Y7^7[cGARQ,VL=KW_M9E?Q_I=>N9:H8PX31\IOQZ)4#K#AWK
KDHcNZfNB(Ff537>Q^<.)01]CW.EY-6G4I3D7;^+B#g_3ff_3M+(O\G9?CTLef5#
5\+UF/KBU5G,cNR8DXeV;]7bB+^Z+R7;a-8ba/AK/+N#9]b1_5HKJP=/_416Z2Cg
2RHECVP__JP3@SY<K.TN@(-R^=RK;bNH]<cZ@RI\-/fVIZ4^MB+d&=a+8aW,7#;=
X7B+-Xa[PPWSO)##?H2g;B-KB,T3a+Y?3R=]_b;9W-KA]X?.Q+XWQWYGa]V.c>ZR
,f\=_Vd=0#?)V=2R]e=4?^9I.ONJ#Y+GZWRb.)Ua?@JBJTV;6=9MR=g9Q5WT4=BM
).AQ2NLARLQ#G6U1cSDSJH<W]Bf-&Y=a4[@Q^@@O(3;ZSQ2K5J=-b(PC-(KA3DJ[
:3\BbLU_6Y^eYY30\L9dDM1F?;g:P,Vd(/6V-?Wb,=&UagN[MX7;c]e/e3a4FdJJ
9b+:&-+(0TXQ,^0PX@;6MG9=cRB?6f:UT]A25EfS@PB\3=T<Wf,.5R]]e5HMR@\.
00HXVY#8/E^?Pf1]N86L,C]9[PNS2[9^>7G8#+6UQM\(^NJ0DF;/G#2JIWc8ZE@+
7G_?#<4)V=GG=^bQFG0dIdDA&X25aJ:QdHHJM<#XZ(b?cL/=4T)U3];Xe1>VO/<Y
9K;OI8b,Rc8\WRYc/.DTL(c,+g#T[K#35@]eYSf(VJ,\8LOZ:R-P=FDX.aL+6T2Q
(Z.N6D19Je/5E?OQ0A-UUQEeS]TJGT5FFb=RNUNJ2Z.[0>SLPY-(:GW[Q-N4a@Zb
NPC0[O9Hb<_fYS;:#.QDaS7V)<:#B\+)=BGD[K7\^KQHC@>e:d-gBB?C_[SUIYCJ
=9?8P-=<ce;9X>U?XPP[NU/6@__G(-D&\#\bULG55VAO+1J)YT5:6,;Y_?B7D-0P
0B,QG?C4/bQM+:,EJ1/f-[Z>YOeTA\&>5RSLY:M?:P(d]8^VVe0feaCS14C\R-eD
Qe^c>SDB^FN;E85B_(@g6a/AGNWS05+Y61De:We=C.#HIYRbW3LF/aQ7dS.=:3#2
]fLcDZMMJ5aW2b9aC7C@aH.U7D-eUVHBJbIE=KFcL=.DBcGAY8<S:a&cIEZX8LBI
/3+>@RObdW;#)H6Ad2N1?HI0daJH@W-H@_(8\4OgdbgQ/;T41603;HQR8fA/H>3@
1U(#P)2T1c3&Vf;=7E;R30D6?Dd;-QgDFTU??06d6[JY:U9J)XPBfHDEVD]c&W:)
]\8(,&cA<eRd_8,_V_KN6Q5>SA[TF&)(E?0:)8>AV863cbDP]-8:7V:[KTdI:DKG
;^=?-]U,D1=.U;gX?\@W5[3ZR8HZ7I3E3OTME1>]#KV9KeL-IKd-Y^=\APM/d&dg
0H9X5fR.W=94U2#H]Q(dT:QQA(fGMFK\0)/Lc(EYP>>a348-<E2T+MNFSUS9DS2=
9&P1;_2XR,cP.S-^dKBV0^LIZc-fDSXc+N8fc5dSD?[HGfKcSFRIfW1U7E^\+N4L
:Q<M0XU1)0<&JW:J[-2[H&[J0M.6.TJ+g&D^GG]ZT=AE_#N6.:9+d#LJbZNQ?K#M
6??f>Wf8ZOFCdCP3GJ9;,:8:0R.O?2^.6deG1WMF-]f8W8N#@[#GeR4B@aE9KMFB
]D;9=_0H+Bc;4B.DMDJ)>&QHI6[UJ=83/W^/<S-bYG^8&_\a908<DV(ME2SB@^eU
O\?V;R<;cHd&)=[He2G[ce^QJ;8eRZCZWbW?&OYX;^Cca?0KUIASKVH+]FWTD6^,
-SN1FFH.fT4072T1?[?QP&R#F,P),R(UTF:dNOQM4J95C8(N</6?#W7RG=Egf/PE
abMQLQfBC&c&?2N\J.(#bO[d&W+VWP[>]Ec&NdPG?P<R-ZGX>#=09=6L;?:(B/6f
C./J8E89H#c#<OGH:P0TBe:.N7BL)HF)eaUSHMe#ARfCG9gWL2-XV.L]JH_CbC]-
L89g;&a4GHgSHYQ;fODQS_AS0SdDGR7GYS9U3G+.d:GO#,NG4SV&&&].F9UdH_YD
>5\&/M)T@;^Kaf2J5ZPQ=@f=;S[]0[TbbXGHT<>#gL[YIZ9f/bIB[?05:/?RI>UU
YYPg&AW3g_\+gR&M@3^cLI##d9R[3aZ3,>Q=&d>CYG]c(<f/A,,@S]5P4CYG>5:A
6Y0VHb(Q1B1,E1;_DK]dgCGR]XA3/H\YC\Y1aX=GHb(a\G?\#QPUTHCS@.F?MZTC
#G#XJ0GXg:af2P^?;F]ZUJ[a&-:B]Ef3A).c)90,NN57X=KJeTLgY6AJ8>d1,G)I
a6SgK2fEH/)ac(,H)PY@Pf)IQC>GIcdR8Z6X\W\29EXcdVR>7c^75L9aED=]3U8H
_LD]<cc\e=0Y[9OZYE^:6<,NZ;C19e3c]_2HUB8MLc#XLL0+/Z[=TUJaGV>dJe\1
G9NGXN/Y6ZD,2cW)HEDX?30GR1LQL#[d<^Z@+5+Se>6),D(\P8S#4H6O96+cU1f^
&Y.gF=\HT,?82LDO]3T-Y^-+PIZ[dB\25&/f5[6C8&UQRY3.GM@b]WWg/Z^C&c#H
PD,#Y48-/06);WfW1WQ).bLQ+@)-/W8D5bbKQ^g[5YV[#[faLU#M;J[75ME?Q>6M
JZ5VX+,\G6E?WGX+9d_M44L&GNEEY7Zg0^ZH\[DFE-e;_0B\OU6WJ,9+60T\0<bU
O?e+,2R(9YU8;\<-KT4#-6)&R_RL)61)e\NE#+B=FPR[@X?[:<JU6M9#)P?eNXO-
[4[(T)U4_841e4dF[Xg]a&2W#=AbcN+>\^eg8_4?P4._R,;/V7/DdQ/a.XOF>Pd0
-)F-+dUaKP\/dB@QLX\W02TNKN^F?&,#PS24Y#;-N7#_eP^\PU:K1\O(X9;NZ>@Z
8EG580(H7+gI#9\5NC./)&J.HWS5a)B6)]g;<O/1(a\Q9B,d-:T]2&^a+7FBW)/W
=)I;6LC,_/90dIQC99S&aK7WL.4LI^:]CXdHO#01WI?3dHa+MH/]K[f4,SPFO[OT
6IbWG<dRA=dEd:Ba9dWd0MC[Y7?:c:(?G9#f22,U/N(.@<T&L/XSTNK0ET6L[J(+
D<J5&\>HH9P:#R>T1^cRb;=[:Ugc_-d:S?EG6^&V<)FG;W^:=F]Y(,)2a-,E/G?4
07aCV:PFC:/)1fMGgLH+NM?N6-XYSCBZZ,;c.aRMg(M6S9YIXY<UZ/K1/J(Y@N)c
-:@_#];Q(d3d4)#6Va:KKJX-g(<5a/V8=Q\d\VM/;MeG;@?9W4AYX#SZM&4J4f+-
?XD<:N3Z_1L/S??1+31SU)CRD6;G(C4+V,R#]L>POOKDDW@H@-Rb^68Q\Md(GR3W
g/:LGP23>#fSaZ10I_RaeRec95T5X,_@J(6?A]O&[5^B1Z\US:(H;D5PJRE_Hff#
DGHFHBO0>FfgVH8-IRZDcgPR?]CQU\:4(JLQE4MZ^4#MOXNE9P6LdaR\.Qf;ITKP
H(7X.fT&M0;W](g<]@F91X75RHH?<O)&.SH3)7WYFM,&E)&aZf5=L?0JX;P+JZbJ
_:W6_=6QODdf9eO7UY#C<<5=_-LNJ>/\IVJCEJ,AZR9EX?b27#BHX@LL\4FD24.7
@^KS)F8fdA0)#YPJ>RR9(ZNA,R8JWF^I>X]W;DW_Pg<c2f<V#4LYR_U5/c-UQ.63
<]HNLA_:16&W?5=d(T=Cb2XKBJXeI-[Q^#=1Mf/d5fS[]9[CUf8,N+b0O&Ad8Q;c
:gGJXDc)=/P6_gPHV^Z)_T]aG+.AX1K=185VZ4cY63Q<BS+cE,&SQW\K>H,KCeI)
1IUISb>X7RV9V-dc1[ZPUYE=4+Nd,_E(2GaM5?@OC<R/&SADf#.<d\SX0G&29?KW
+8EH5B:F_FYf8>PO>/^Q.a2C#VF2HN8<7?[#M,faU7?GgM2KD0_:I9?][C;8e&>C
6>IQ-f?_fBE9KS(&;Q<RZZSVafH0#8H<bL19.Od5S.(C>Z>NBOD8?)\fa-453?:P
N:539V_-.1^U<Fb<[cZ.]5HY9T()6aR)>1cJI8b8#?3;KdKQX)3QGOT2c]2eaV1_
Sf=Af9-Q>1SU&2fYQ&G>9A4CS(e,43P;2g8Z3CaH8NB5KXe.TUVfBc\=eO7F-ZgD
.V/O#W0eGRaT=Q6B8-,U9B[B:D(6ZX;_@TdUK4-/Ebc&(CL3I[<.8J_&fFgJ]JJE
X6_)JaD7VNA9-NVOO]3=_1N/TLF#<,KPXI.;^+b4b9>\^<^Q?#@-<C0Jb)EYZ7E/
A1JY2.E6Q=QQS\4Y2-HI4L-^MX)83WY6-TGU1H(-H-5MGFRL9J0._R=]0SR^cHb^
;J>\=2;,CD(I5WQ-T^GH&>M5:ELBe(Q:PG7_-XDb.ALL+@9E9bWL4W\X)2MSTR@C
4d6^81-GaY9Ig(3UC(D[gUM#dW,(VFERaNQ87B@Ub#6TV=BMYJR/<4(7N7KQS0KL
(0N=AH6ZV7&0Z70DCe2OSg:b<#>b/ISb&D8(#;([C83^0GT_\4_WKS@_C?=MO3D-
7R1&Jg-8?Q/9c0OAWTAbOX.#Pd9L5V2_SZUTa#0dPX[G\+b7753&</@I97e&+_Y.
/#:Eb=DSDKb@JD<I\:F-+H;=73&:>72@=Q4VO#02/.\A&JTPN/8SA.X:Y3<O-#_V
]c7-8g:UU+#Z23YDKa/BR0RZC_3C8HV0Y)_:Nbd.CPWAK7:Sd,?+#MLUIV01CST@
=\eOeOGHaANF^8--=cOE=9#3X9F#)Q\/G22VJDGe3<V_A@=1(UM^Y.CKPc38G>Bd
KJ=O8)JM;;7N]F1:dC034:X0\9FfT9-f<U4<;-&.&=b1/_ZC^)@H?NSV,FV/[N0(
cCRD_f[77-32W@ODFMT6L5\RZRV?BU6C3^S9d@:>Xd-1@6PDP8#I_D^\a7NZPAd_
O4\73GCAV2W^V<?5\QF11Z/\8,#\I?NZ09+GEO_>TQT/\\+\>;5/C=[IJ_g,@(f&
HD?WX?Wg?TV>=#ZBU\(QZfgA-Wd;_TS)9cJ6_aeN<#7M0+]Vg7GPS@/5BRf\UBZ-
23\YK^g\FH(;&KI?KJDUS,]S9MSQ2fQFPc@YCNWBcC(8^1]Hc^aKgH]TK\WO(VV;
7K_bE#FU3K)^)4F)NgT0VVSSMDO]9VU@ZPdJa5DJ).M\PNYId6?Dd/g#P8bN5/2Y
ZIE86-R,84UP(5TBBVDD@.0U(U7PY4^Od?8bcSgNO@N:)bRaZB^,UN2<LCZ(+(1^
5b._f;4Q(7PHEBXH)LE_7a=7IPbKd>T((,&SJ.@dE/(>a,I(K6:M>=.MO<A,d];)
EJVQIYAY#3d<BHM?)JHW.[LYLU+D3BK;fVf3;57EfcG>Q#a[G0CU[K\&UZT4?WF[
OJUXb+IW1Q8?S7R/5;D[3L8<4g//=6M0P&KLVY1MNf+3/,8EZFgZJF-]0DWfL_7a
RcaX_AA+;>ZQ_W.]+QSN?UL&;g7-]g;>S(S5NCf9CR.<OYR68I\E:8.W20L82+g.
D[H^J<A9F0/)31W/\W1?&FZXVUI:S&:K;9LX+d5H&VW[g:4aKQ+RbecOV)AK68K;
8UJ/TN=:04<UX;gDg2S>8<bScXKG]dSe?-W23H&&X;6=@51E-B7:-.AYJAE7+gb+
Ub@3Q-^XS#&_8)C)_WEV+E9I-+R_T[:<TP<RM(_WXM_R=YZ//T@d6=7g&C^F?SJ@
F+TEB4DXU^1aF9cHGXGZ(=-2-ZB^aRTYZKA8>00=PP2;9(Fd^L0Ae@=A8J2JTS0K
V99PEP7?@.68Cd([?;B_^SC?SI^7+PSCBTGLEI_g2?L@]GN2P&:GUF[Ba3I9dYa/
C3@M.R;gQ<>#3/U?XMebHI7e;DZXJ&R-N1Zc.BVNEWYBSYD&V&&6T7IGf)H/+gGG
WL->B(T]A\)aR+RHY1fNG4F>5RYI@g?&^@D)Je??V\9D^QT_4GO3LHd/):PBb1[>
^YM5@N:3D1Z/F1D+deP+F@[4-SeLCU>XAD1-^WDH8UZ8F;bHMEX\DO=dX]9C)b))
4^OF&;9_-6EA7CA206^VKKH\b0LI1T#T/T/;_Q63K;N4C+/g(T<29?#DI1a)-[a\
S;6FI/\[,fg[fTB[N?D(/8/-E:Q;FJbbG7V]_I0#_24UJ,T^e.L#c45A4<TW[F+8
\3d&52^^.).dPI,CB3ePGCXeD)]:)W)c\U@\0e2]I+f_6e=.^DZ_c1B7\c,^[@NJ
5c_dC>3P&3.baLFL60@7J=6BGI^P(4e30b73)cM?PMT-<F)9bcW5&Se,+g;4gUN8
eN2QF=],Ag4[&K.6LM7O>#JX2-?<Z\[NaNW2WGHgA&#c+S.@\-8TG6cQY2B6=ZR^
=Re&;e2e]]N,O.YOB7_JA39X0e[3)GFLR#W)BC+W8,#^OMBI@2MF<K]Oe+e&bJ#?
Ta.6IZ\M129Q=4a5eDaD8FM5AMfEM9=(Rc)<;U>C<QOZE<CGCa:W4;6TAQ3+aCG+
IGb;bNf/X<]>T4[?70GP.B]&_4AT@[B;^_:M9XJ)@)8\2^3A3f<-BDfO6?IBb;]?
2LSG#DVO8F=<[AfGUcHF6,C_\/#b[?,5<3JQEg>,TWP[4O4O70=4B@OZ-O(OHMCJ
93_YSW-]QCSF::IFH^@]VGLY5&dSQFI?K)NA15c]NDQgA&Q#c[7>/=Ff<>I(ZTY[
g=A?79@JaH+J;)#U.2UQY0Q^f<>BY91MeJ&^f(;9b_\f.bK#4@:A^@\U;Of]Id:d
2WFB+KTE@?&.GSB(.A:K(@fF)&6\?>Lc\?P5DTLCD.1?8>+-^V@PVee@-TA.[f5U
;:-2GQO2CC[MAJ1S<-K\CP,#bG,9<a-H342&Nb<__VIBX<58a)X,ca]eZW[.E_EK
QddTXWeT^+3HBLM,CA<g\\<EUc>a&\RJC4g=UFETIfN7?U6BC6:YWWC-FZ.4ML>)
41)EG+LfHa(SPPY3-V&](0VPb?FBYbKf/R)#.R&6Y1T1GPb;1W6W+N^Z89J)&,)I
9V]4.EaJN-8A5ZU)+(g67V;?2)LZ2J05@M,&>M#.J>b@:M9OKCR(3gJDNa8.edM]
S&L?ZYQX8eY4)RD6C9/Ug<\@+d+R]GAU9d^6RA0G<O;e-2VH,Z[L6(W)N.A:R^9d
1C1G(]#IAVJ@V/Fa&#L9)b5L8&51[-f4T_P7[=_PIVZPbXHdJ_[:R4e\@3W@K?4)
[BZfRd_18^[IQ:XGVL;aYWKP4-IO[MDB??aWeQ4(NXLa4KFY>3HGI/eC9S);@XeM
3)8EPg?BZ6D1/H08/E?@<6VI:O[<1B-#d9BYJ,2B#b9(Q7K6^AV=>)#QE\RJCM@[
HFG>IFfg87_\?9TA0\N-O_g@=6c0?7)Y_5@6J\.N-^D;dX3D\E5gdD+^9X3F#;@P
])-3W7?gA&YE;X3=WYLB(<3SUM^-<_;G3Nae2SNN_G=4T_36a#0VI@bN;5cO,SFd
O-HJH5fJTVdCE1WGP:dC]3\DTM9S:(F.4dELg4>?)?3JL[XG.T9?WIa813#H>I@6
1K,F?[[f<I&@Z/@T@#8XK9)DKJSSZ]0)>TB>1MT(V_?O)@aQSH::LC],84NOe_F&
R5-HfGE;7-[gB[N^dT<37UWH@68TZK=ZFEe@4==86)V5b7W9aUCbOIWX3Q_M3HSY
LTdX,^dF3-AIDRDf(--XGKCdJ7/;XITdAV]=ITT\X&?I4@?f1SF.g?:eSQ8-]N;4
AL,XQD^:cR<=W/egX>;]GA+_Z+(:J+NQeQI(ce(A9S00Z]g#b]1.7I[d>-O,UX)g
NG)GCYd,^=F9[O1MR)<I.>A7+].7^\?:T-P^g/@Z2:N9+ARS.;DBIS10?7]CU=CR
=)3^#fM4Y.=?IIXcgCP:,ZTTI7>\[P;Y++F4;K=g+:IMY3I/U,&\.JB0WcADXAA-
EA[3X[F_QDXS_^N:9GG2U9&GX:9)97(#V]_8;.O_cd+<6I5C^,^3R;3U72)T?b(8
C+F-.CV_7A]@>N-TPRW==?IIB-+5,]L>D<1f,A6Q-HgbX&:S+@K3P0;ZOMYHVV.E
B&E:3Hf4KE/\7J+b9EDNAg)+SH)C3L:IIeZBg_X-6PH9?QQ,]G&BT#]UG_VL[&PX
Y_\a^M8cb;da6K:_B;NT+VH07d-&)(YW<)638)AAO<B(8?=X+^JY#F3^[fII-5gH
VR7gXF(3&T2RA+c=>?2W]Q^V?#M.+(@f_DO]>1^HgNU&X5@QDFb7W2C5@7ER_NDI
;(>MY3R0I\SW#)Qc[(P8Nf@T(gO#=>/A8(.M/WWbHQ(c.639-XO,,YbGfP&^3TS=
G-EGa.RX(2a[>\I[5L?S5.B<f/Ca@:LB3c(@9VGV_#U.2eQ8^R(\)]4O0F>NVH#)
#MI38(IVRCVc]TL4T8-+Ef_ASYd(2=?eO+&3CSY]3>[;9.O[S?4.YBE[RTVP)7T+
/=@[KDg4<9&#2QXJ_D<M(K@G4?&Q]Dg[gT?H1?E[V[B&..dH[0eP@Z4@2=V5U9#B
,&GbLaKdeY;HCTIOH59EBC5_E3^,48fURH0E4VTIT@>cGa@#3PK)R12^G4GE;EdA
10]L9?N>PS7OBW^Q<dIELWQWFU&=&]?eT?E8.5>9(LXS)ZLZB=TX7ALI-WC,<RB?
NTO9<6J3)Ydbg6,?bR9Y[H7B>54BTHM[XTD]U09<T,,B:SBcUX@\8&DW-Za\XDbg
@^0?Tc)^7>.FbPK-P>7UEX0#Z[L>gRH1U4]KK+c,7C\\0ef[;.3X.d>1;<>/)NY\
-FG49R8(?>=aO[0Y]XA3_)I+:CbKZ97#,BWZ9R)(F-5&KO@OB5b7Q@)[U8XTX]:<
M1D5#,[B92:9,2,/IPLOFSHO4->.&K[-VH\1PU[GI&^[aI<,3P+1.Q6CVXRJC4WF
8?ZVIT),M6;J])&Z0X157VgDANec^fL#F2F[D=/J][5V]M_4GFfdB3ID<NE6][XT
7LL>fc9YSG:T[8.<OdSY;+?GOe8C=XKY@b3]VZcTTDCV@4>gAF20,4c(-W1EYbLE
?CLB+4g&MAP<KL0Pd+I#M>cg\][TNO2V,3(L;N+9U8<2a9F7?:L<WBI-PK)bT]f)
_a#8Fe8aFdU2F5W#N>D6.OZ5_f_6],O_YS]DGXe5d/@?IL@&S(5Z#4BGM.AF1Qg1
DN1-#]\O5-0Y[7LX.f+J@WQT1705Z)]XC2EA9Q^5f\d?a296EeZ9]LREd(PKBV4O
5>9DLOaM0J]@Z7-I:AY7(aA8eR5]TLE,K/C4JT)DMPb-J[f)G:]+g?WSSJV>c?9.
Ta2W1-)aRc-08;?X(,TD<.DID1(QS>Hb^2]B)J26AI3L[:?g(e:2NA]A\O>3LH)A
_3A#AeRN^&[5SbI/>UGc/e\af-K]fG?<0eGFM&/0S6X[L872K,3P?=QZQ4-SZ(:7
B1df0Q@0>._UMRYBg582EJ.2L5W;VVY>GBRKHPRS=\+a^8F/3@Nd2ZR9e)g_SB\9
:H3-eU0#0>#2cSc_8#4DL8.4>(H?Z=(G,K1X\T7DE(U6J7[^e+:+&5,4V3gBaK(S
1U;8_,Fe</^D[bKCaFP?@7I(ITY>OTF6-IZ=5WY1SS\/+C@B_UPc(62@BIA-EH15
T+G2Pf05K=SZdXbH_<5(8H)?_\TT.<=FC(fCXUL>NdB7R_4^&)BdEL[Kb4C^.ed:
,V[Y2+9+^C_+R=e[Z)U9]BO<U0JO1?#bC[>0/27-1>&.0)/&2OT\A4D3Qd+DXbLC
S=:IfI#F_K-(PJU@[aH:cK<H/CQ4H49HN(#IE7XG5ZOb1G&;AS>^\L4SOB&YOTBJ
3^_>+64f@66K,:;&a<>acd&V(S3PV,aOcHE\>Y>F\:;4TPH9@8)DQMCUF0g(7d:=
X^WG_:D0.GGHb1.3QFf;)e+IbfS7XPEc/\2Za+]#f=\@:7aW#a.;7=WF5]W4Y5LE
D#5GPQCgJBTVQ99(XeN81-^]<1[8>R\Q;[Q(M7YL3>:Wg#AbV#c6;[5cUS=.I#?f
;\3aYB#C1.eUMC7FGQW^;JQf.CRO9IF7QN,D)aR+(=_AW(4Qe,BGg45N7H[O2HFd
/ND=KV38:E11_21G_VK3NXCb4g>+7KESG9=35e]7VNB5(RdJO9#?0E7cUKC/^J97
Jc]7W4S]/;R]C8:dBc7BO//SL^cfR;BIO^Aca/,=>/X\-+FV)KI:)<R0L7Q(d0HG
?(aF7YU#Ad<b6ZHa3=H(-9RB;6<GPdED?A[SPO?[8\A-\1><=?FW[8YeI.68A5dB
L<2V35>A85<]&J,&,]JP+Z5e^..9ZJOG(28AD-a]7F9?JG0>HR4K?]B8X\AET3EV
+W.@:f(\P@SB)XJ-AW1a9)X+-K53/bdZM(+gGTATRa5<2F:V[O2HWM57]g1.W@60
2C-7f\B8.cS[-C^I9(<]TMS4eMP16>71YVYLQe.K/_/g&3?cP2Q0:YZ-PMTKZ+H(
P><#OZgYFV-+B2f=&,3<O]eA)W;\3]aXD0S^XZ6SOVCO+BH.Z+:bZ;.)(0^@U::<
._N<d>.g09NWRQ?QTa]YH4:=C=H_\C\H;]U8#1W2d1X3[eQM;f]aK:.-JF-F0IM<
8f^YX^_8LgSBTMGVZ_[d_Jcb;ZD1\9a+\DIVCcM0Gg?;+K[</,I#XbcfTbfIW9QG
^FB3Fg])A_Yb8M_^S)dF:5>4/L2fD#(S72>L\IF=)]4ba?a1N]?gZ,eIJY(J/\3O
84Wa]MA]._/@Te#V668LBd9gI/S1Z8PcbM9BNO=H-g9,M/BaWE&C@U&HYF/#R/f#
T8[_G4Z^dgES<Z^N:Ic,dX7gX6EDaILKNaZNIg0=HMD4\VSPIR48CBO_^N>;Q5PS
E6)Kc9+)2Eg&5TLV<aGf;4,4][NS==D1P1>H&b]_UfPY7\:b68BNcOfGR=?N(0SX
L:0.J)BPFPH)8fIcA[A_:c5^MX8;aTGG\RKN6^O6]eZT9.@(KN&\,7Md4d==QFB:
-fcZFD>MUg7C<E1g;AA<+^IW>aW(Ib6_d4PNU.>15_6IH3X^])d-@a95e-eSe(1>
>>SH_.d0FVG1RCRCBbSKgH@7.7UKS(g(cXB0a\YdQK?C:W<b/^-Fa&;-^Z?NS5S5
\]M@XE]_M:2C7MM+B-RQ;f=:5BIJN((L1B-Ia:<)0ZAg/H^?KdQ6,XCCcDF6Y\b;
f@aAfd/AFT#OR.=b8Q&2-N:YUCL5;I-O(UJ?fXJ\9:3^8d]0M/2<I>S2aMN:d()g
Q^G,6/:R-NP^c=ZQYCW@f;KRMD0&A5PAZ+W.ga^KX+U&B^Z<a+aPA-I<e7-V/QAI
e#,LSa64YU:>D[Y95=WY2V<&B>^;ba9+R#_D,C+gJ8S:<M.PSc+Q>/>2WKM.XTfZ
283^f9^gXI3WFSLe.G3L+ZF=8Q(bJF7H:ATIOSO[^27[47Q?.CE2;32;KS(>:>gG
efGfLQYP\>86(7JC/W?^]-ANNQO8+9;L&)Q5O+-F0Z/f8bG=;T=(46-eb4A[_MVf
[1C4)?Z@WOUNg^/@Cged0@UP+4WPV,VV)O8G\C/4\@\MX8SC380[HDEKP>F=@I]O
&HU\=(5CBa+e:,[3F]96BZX?)+NK281H:+M\]beP?R)MPF,\?MI29QE#g9HbP84E
E)c8b8]M^RcCeZHFOd#R0Pb3HY1)UAR_TOLGc+<]ae/3fKDM7=dX.UPESBL:1@aP
I>C+L^&V^Q.PUNcUc5&=(^.HZTCDX,-)GC5L\</QWQZ6<W)[3>7?b.DOFRC(V?]T
8+gUT\6[DfV+g9G;N9E39&0Y2^OO]H.-f/SEd7ZM40b.=CL]+3d-(A4(Rc\e:.eK
XRAd<ba\_RV,#,Q.JWA(=Cd)SK#N(d@0RTF/fV5T4;R]<ag^>?@UXbRCPR7,<UB/
3TAIb:_]eU^R1-AbH2IBGHWZd/FaPD]8E&;.H@[N(fCG\g/L0S7E2\_M[_M0D(,/
HH5)O\1#GN#R2_SFKA;[5f4EMK&]bP-]cJX+(g0D6]_9^35PJ8CP;&4A&=9F32(X
A+g^[^UJ,Tc>T?LWBUS)?6g=F)>eB@>YLM<\S30,Nd-@V3gN><8(LQ>H=O5?7-eX
GH@d(ELA7A0Pd&7K>a?@P[@a:N->A0.R#Q#bH?DRPBYZ#X#ccZAKG+^B&aNW#&^=
4MSJA4f,0X@3=8M[\ATfZ<.K1>0#TVKe/06E_ba/>TfB:dfbJE-L-c>OJ(79OU[X
1]YTKONJ_He094U[)W68SSM[Pb+;7)PEDaX5-PR?RATa,0M5QY7L^WJ3Agc)CFO.
2<24:M:>f:??a6_(>eNI=#&(IRW>7[O15>+,F9A-H,9<?:bUd&>;QbEDU.?1g_ZO
6CRLSB__>/7<44Y=[]H??NO:aQJNZ=-(N98V#;AXRX:U?:1?87A-:aTgA.SH_[gZ
&MR8>E8=cHLf1P]7;/fEYTK8c^;.P:c[S@>)1.I&RdDb]gBf)33@(cK(<5CaDa=:
WW&:7?(CH.:dK/=NgOSE;B^Nb+g[[Y?Uf7:Fb+;Y&H#X<^+eG@8U_6/Y_1bM#Qca
9V^<bHcZA.2-7gS7b.3K]=WG8#O8?@;6]_LE,-UMT)fb\SK2?]/&U7<RZTB;R=27
E@f:>_DG3P;QS@IP7722DbM-S4:1Ze_2+(c8YE30?NNH.7H25bRGe:<[4PT8/<^#
3\EV#c.B)]g<4JDcB1:K:@ZfB/[OWUWCdA]A,JR,]R.g[-e8;,f(fb&OEg1,GTF4
VA(O/&e#0XM9YJW/BMfc4e_+@f>aHFDR1_3^2=;bY3MOQJ-GW8e1W;S#[\G3X8\_
83TbZ<:O.?OA7<9+DM@[([,\:8eS1Z=S]A>N+-_XbJIJLUB<bDU0Q81]&NL&1aIE
54>QXGgSL[DXLTK^#9AA[)f#aRHKdO1&a]WV9)]&9b,+OH\2O#]M0]cbR:GK2_K;
b5#>OO0T+_@9\#P;0eeK&@971YI\1T;<JB&Be0922dH6a4Zb/f9M-+TEAQAeBMb.
&a:#PRL(X.\bgL,^_HT(JJ(I&W0DdC0D<RI.9LP3IU:\VGVa.^CJA95c8#W+J=[U
62925149TG/38e5=2Y/H2T/<>DH1YZ38:cSOG0I5A]:6)K^W4124R[=VdcJUb[:?
V^B]SBZ?Oe,65bP<6Y6Ug+(H(9Qfe@;(_(SMdC7@6I<e2E&L3ABY)F.PBD&\>.G7
CS\8>e#EA1ZcA1@(3QG:#J]BaS#Ea7cgEB4IWgH/TEQD]eA+5\X.Y<>TKb5?]]@(
,25:#E:]-H;)0:@^&]HGNJ1B7SQ7dZO1PJ#GW:D3P]V.@A==T)K67-C<_P&g<>LE
KJO=F1[HMV>Ff(#HN6b,]#EdDIY3?a9JY5d,4L99@DX.d,SY(=B/ZW230P9>>TWe
PDfDf^]--FJ6:gI,T+G&d9T:4L<=^=2(DS5ZTdBN;1Q^?eDbDFE+^@5T?G?Y.UI[
SR(8][6\J\4^L?AK2-.NEO.Q\A;(Wa3YdB+cK[QLV;#e(MV3YSNU-4d17;.ZL_Jg
<?)KZ,;UgSd;13=R)LMX4.@310Vd^YUEGdGQ@<;2eMYMI//D-P6.a#B5@C,(:0)9
((@B;9+DYB5:,:bI:d@TY74-fKGF;RFIQ+.5?\efF\8T9P?0^=X#TaHL3E)(5IOX
?X-)1>[GO+gJQL5c,0)B:Ya(+2TV1AgDMF(J?Z_ZdZ,BMLb#K860.WN9GGG&DKWW
E\G#<4Q?3I1Q6FBf2LB\DY</GF]gK5\6d\0(EB8)PJTS4.;,-0Q-D\,O+EBC&a8D
E1E(bg^G5HM)//MA^d_)4CZHBV3ed,6O[HMdQ3GPRA@fA6\DSaC^?8B<fY,;[6XG
:I?:YcQ7DW(H6?Y:JCSDf,RI>Td(9,\e<9P=@LQLI6K@PO9?M@QdSc37_6e1/PHB
KF]9<^-Dbe]\\\66G:Z=QcGP5/0fAF01>C[M,0T)&E:YffC2D09;EQ.2EDIW@^Z0
G/54eLCc<^SCKO^;ZZH179I9K323,B+Yf,6F?_3Ed/,RGG3]RI<0.^f)a:K-ZPMb
NVG-_4Aa_E4Z+dHc3#Y\?9#?841_^;XOTS5O<b7C\](@#H)BX(YcW[6ZQAUL.\/;
1aTSUJg8&Ee,J?2LbFJ<=a27&bOXeRP?.GHbR#A178LL6/A93KK2LA]8&JS9A.NE
#:J)DVENJ:c-ZKH.Ve(9TKS>9FPc63c143)WPOV@+?0V&9WIP0Y#17QW(?T9QCD7
=T-^UO:DB5#D<aaJT/7FU)O>,DI1e+=aS:ff4)_B1FP(>&T:4(4?85Cea2(WMP+5
K)@eXREX97SO+Be]EXSf2WG&E2ETbO)S-;2]N4A:,EE<SJEE.7eaf(e^OOSd+/4O
Vc^<D03dY+<O?.>2U2V-TAV+S#O9;VJF9dNY>.M88]+U4-S)H+JT:dT_T#[O_fY3
K+c23,&82,<Se)M3UE<WMWL4P^4a=/cOWVDdb;M@6Sf[+?d/&c\OVOb8MVJTB8XJ
;U)WUab)H)<3^bf&3c+^)JIfIb75PYMK:S3)Zd792,P\W+S@7.]IA@BOX_7Lb.:4
9ZN:1WJ(c.IYW@cC_:^NHSXeM=6>@T6a7GC,/<VZNULIb=AQ2L38IQ/7FdVKE36G
^/MJYfGG<a39ZH62-F]:N6N)(b_W5<a8OaFP:=8#+Mb]#7P0dL1=Nf50A7^PE6L[
,<gAK.aV67K3G:\2.E+4?EJ)d@IW+DPg1V(e#M\Af+^?11U2_4:J3/bX,3:a^<+Y
Z-Y>V?T=?0X6T0#>QAf1ZA9fJXgX:::dA_^P\MI:2F1@U14XP.(Kg0S.GO?9@^K,
W:VgT\ZC7Rb/20a:FY>7a8_Z@<.KHIWAJDW[13J=ILa(&[VGE_MNLPDaHTXf_X2,
R.;,B\f;(]gfKI[NJWZL:e(_&0@[XTFALQGe:C&.6&aN=YR&:_CY#(/743#FLgJX
:M)McBF961aJcDQN8R7]T=7gI^X(AO[I95)I=IW/Me]4ge(+^B[6/7[YeWD#b/DR
J_:+.0WM]@-61N4DT;YJ=K(Y)=1;KY]1JN>;N2]/8R&K]Obb:dZ+NY]A/;6eRge;
U]YAM?b2O^/JWBcEeAP7CJ/NdcK>BK<R8I<KOUFDV8MY1+a5K\AV;WDO,2&d?7H=
8&WSd(B)ZG\?P@5VF^N?<@DWEga5-a9O0<9MUKad,?SNHdM.-50J?1g1KLg]6d3G
[2Z=E]K-+K87M/_/+<(I\)B,CHBOZbTe]g<(-4J:/Wf\61eR^&XRAVF6CO<Ha@LV
XG]7FTM1=,262WA>8&5db/TAZP[.SGS&N1U&TJN83[831)](-CA5_#,=G+LV&:dS
2^=gKa_R+U,-PW1X^+KWSYZ_KSQ2#DdVB<N_6Zc/4H?,Y+=T:+M/^8P_W;DL2EB9
LT.I8g(9SN6(B;<;9Y[(T0cAPILO1_g_<K1GOE^)@E^&E?GX?b4/0eZ3#0HFHUFO
YDX@=FHXJB_06[WHR.MWW>0GDE^W97.Z3_=^^:I]CeR8@5H92gM3&1W;6+O/a3^(
/+gZ9&N7WL6KI7MS(b<[=6XF_QBNG,Ob57]/DX-RHU47EX<e4Z4S.6LHP:(GIE>J
EU<W&)P;^]2d:VZMYc\,EO#Y.S+1)=Y_5&4.[R^,8W70BY?A8A9\eF)AE12.@a.Z
DS-Y)>09C+51J3[2;I;eCT>8N^OICCFD?\XR10^.?YAN/R?A<S/0SZ,V[?45^-0F
>D\C)U4eSWP5BV\9[6Xa@Me_c7IXVg==CVG5IL-IUX,LA:J@PR\[#LH_C\JcaEUD
0H0()+0b(?L?/LE-9PVdD@;B5@0PKeK37ETKNYRXOTCC9USJST,Q[^>b,N;E@TQK
F+^dEf5H/B-=MM#c-00,P),>UW/ZSA>07>V2E<\d>.^O&AN?9225M,Y=UeX[(/CC
[dJSaad@?))2QU#TXRBbLR6XD2=;ZV?@5Pe\e:@W>NMF>8S[/c>@-/1g:G_aQW5^
\/D&Q^T#5-P?7JX[COYT##HfWdR?HD>Wg5::X#&,cS\O^G&T+PU5Qe58NHK;1.Be
]NV9ZX5EAI-)(\+UNc;DNX\@/Wd[,A+6Q\=XSOZ8Q?F_HfH5_K3+QRCaLV/7E2=K
S:J52&QV,;(Xc&dHH,+N.P[/_CY#+452/:0J/H;]Gg<R2Z<G4LFS);YD3,;&<Y1b
I6=-N_&54I03Ic^f5,f.3ZOE,JMbf)7-^^M]D^&L\8T?]XT2LQ8I7Mc3Z7L.Ze:5
?6/[(0KD,)gHYQ[8@([<WMK1+]Lc]A>bI>+&&/7@VaP]D+H+EP76MX)W0EJX6FZ+
AcSKR_;a91A/D//_c_\NK6\Q+;J@+>K<b9d[.@>18FRT\2-RU_A1GE/5]AS36JV2
:_Q6DC>F9\ac:,YU;3H][^TfYQ2ZF/;7L6<:NUJ+[cdf_]TNY#8aI\D/9,+F80-<
N[Md5?-@c&81RUJUBgDYgL\M37=B+DGH=@a>d_A4R2I-<FI,QC/YRPI[0^X]3#R1
aDIa(VW?XH:0<N>DL,eF=O(D3SW1DG-f?bM9]bU=UGQeQVKg;NR2HI&&E]YgYZ(;
gV9.Na-Xe\0SY)-D>eJBHfB7KWCLJff,a.PeP^0X)1I665PR>6Q;>G17E&S_URF>
RQJDQ.K_Qe5PD#g0FNV/^O.CS18f&AeYEV<EJM70WL<&136[,+A0DEc8L+b9/Q]I
^Z0+4<DgU60U]Y+8S(49gD;7gDd@#6=dN7)1OKLYY@I]X(-.L#AHW-@WP,:62P)&
#K4-TRL.SXDY:VGUe&W&b4eAP+76F#.+R^T1f/ACKbB4?-D4&^-YF]Q296TCPB)e
B]7^42U7F9&=4,@>6\UdF;)K\R3E+N=gEcTAF_EKMYLYYee@1dN]ceN34.V1SbDN
0[YT>Uc;R)T6D4V.=J>O0-S]?P7N:C-B5[0Ued3PT(RfcW&CSG<-@)0+YISFJZ7\
4XC(Vb1#\FFFfE(Bb><bYLGHbggD;CJN_WPOgB-fNJQN<UL@d<N#XWRJ@Q+N;4.:
C[YOY2_^e-X4)MHbQ6[.>2<:-@Ig/cg-+O^Q9QWU/ZfZNK;U.PUR-@/L15+U44E>
S?dFK5C(CT/DJC:>Y]^1;29B.a9(1@e#9XGYT2>2VLa)]Y5c5deCUT.<)EM8,&#+
@KV(Q24];+Q4\L,G,2G)9UHC:L)1&.FZ?&X,MX[0907N?<QdQF1[>:+7B?g/+09K
)(V8I/.,#f7)])X\G<\_/RHFa8I3B.aMFM+CI1_dAV/;?4d>_.2C<d96^G;@5f(a
d\R1&O4Va]3PMYgbB#=KQ5ZD,Zb.T;0b+Va<gOM5Z(E8T#dM\fLBMIb4gQV>8e/+
cUKLD7,#bBVYU/>/Q6J+@TM+dTQ(^0EV^MLX.=U<ade#Y)QB7VLK.V)M.eTaWf4]
PWCOD<PJ83fNKCgS]&eRggc2fE)4>VD@d4;>d\&gQP8ZB_U5#GV;W4#D92Q]gfW2
@8<VH?c)OD6)<gb(:3[HXMR\]I1aM,Q0O/@H+L]_5/]K.>1MC>E&YLcc,WH?9g\0
(>94&3&7/;Ea<X.Ia1@&S[cI#f]Dd?\1GKV2N&2&><f+N&871?9FAT7\6Y71+K5@
17BEG&/=cO:fES1VHf+\aF7R8-D+T=Ra+Z#G34NbP>V_-/9\@:/8VQe.]e1<?b#\
=eZ5)J(6#@QG\&e<#><RCeB&4N_#H.46EI&FH+fX>M4:20H5;4=I1[<I+PA4TK:_
L#e5YF,KJ:=@?_=)-<)O.+e9Ob0e#C8F]+.O-Y4@eQ+9.>CQ\ec9b#C=TFUbHVgG
_2HNSG.G@ZG34gJZ4LPKT4F5+YFW3:0-0EfTd7UG8P15CgHN_9PfQ->A3,=g_?&F
;:#1\=T4Z-HT04YWH9@PS:a)R=V@M]=S)W6:[#6V<6R7/2#P\Q<[>\JbdOcde)T:
Z<\3dI)dN?T@B^EaJOL:?636Z[aZ0SX6WH2HVFf6Pc&90(THUa6K/V6OK<@gG-&S
+Ig[76FNGS.>F3G:-\AF7e7HgT;:E=JLbg\VAV6b\,5cY<FBQ\YA^O6PU(FG-TP3
J^=(AI.dEF_g32&+0-FS7FIL3?68N-&bQ:Y2,e=)8@LY0YHc4)#Z-&A<ZM#-eZ,;
0QS8<)[M_Gc@XKY7GLe<7Ee)Z\?@G]<(_fWU\-8O7B;_d6=40/A^81BgI=_XfC(5
E=YNP),MP4Y.BR4dWJZ)E<Z7.=XV=.DeF=HLR2aB[K&-SUM?RFeSG)[CcdM>KB8N
3BC8KC:+gK4aWSKF&]UY@^GJIH_Df?\6Xa#b05/J<d<LHF^+ZQVFE#e/#^Y3W&VB
/GGdHLdF0.82I)<;cK\R_3ae]a6U/RQERGV_;)NeGM#CX5;agWDSRX#K&6BgMO8E
)4W;EV:Q=0O-_W:K>+HSZK37,#8LgT6PYZNfK_M#,@\0</IM+WTa->@Gd3AE<6,+
L0C@L(H2PS<(F9V;L;B<fSJN@8<WW)Z>d#^KT=g4DcK#ZMNXA_XGa(;8_R72J^8/
F+,E/0NRb3_=gN]01CP.>dN(8Ig/gD[UFb^;LF@7<NT;PcWY.dB(Gc78XJYb/\E#
4Gd\VZ[@=E9AFZZ9WA)JLgIb]Q@O3+(XS117\F\0XLc4dOG=V>6:(LO1HEc2P/I,
C\O0^XAd@B#^VbPV&X5IZ-07Z>.=#(A0W>d1J5#eN:KTY4_#ZVK1F68#?8e<G8;8
E;c4K8Y66H=S\6XSQW-H3DLX\4A_IOMPgZLO<&Z?c5bW3\UXe5)20ac_Ea24a038
d,5CQ._?S?bf763(NaHRb,[bf?LM_K+&ZV@aH6VTcCaW&^JLJ63fTC=U&#;43A)K
\-X/1I^4UV@^80Mf6Z0^D(=RK-(7KJdI.NUd^M)CZ;=Y?=6_X-aB3M#/KaZ&1V&W
#Z0d<Jd?8;c-)eGJ(\MY\?cP;],)7DDJ/SN)ccX&E.>Y#G:/=d-E-ZfNB=Q9(UD#
)P?\\HaLC0UM:E_=YLBDG0T[,NW;8&>IBAc:DEU]7NM<<C^?IQMIJK2>@/Z^;YT@
)_M,E)Y#g6H]+T7^=F,?7gdTS;&X_[@>_d>A\)a-#b-C1CUL&(fY;46LV[X;G7+D
ID+gfdcbD^Pd),g^1.WT<(J(<3cEY;8,)_>&(\HM&Vf7DAEZcI98)JNO6XAbTdS\
RB&b\J:.W]MAScTg3Ub(SWP897)C,gObT-C:.U+[c>#4c\^@1RR9[.U=K2UG+N(4
Q4C7=XE<D@,TVE+29(HQ>+)GbI0@-<N_cEH-9c>N#Y)?=XV;[c_@2=5/I(:cYE(M
V]O<.g(&789g)Q1U]MLTN(SN;MMKPLd[EQ/OPcXaY?dH<OU;0CUI>W.8&..,>\[_
KVMR//F\?QAdJTL>OKIK;,<NW53)LVb29RK9K\#C3f3_.[Q12:b/I]NBQ:aR&7H0
=<TG)__7HP(6Fb:3><C25TL:XA<^87[a:GId]?Ee&13JZ)4V#?+.eK9F(#F[NUGV
\B6TF(aL#CV9Y(VT^\?CcHD>GY\SMd,aH1U5SIX<X>Z3H[a07K,dJU]5PR?-.CBZ
591(RcLTAR]INW^?66;,FX&F4H1?0,@:1/#Oce2O6ZT2MU?b&)FC0NS[cC+:O<&]
B&[L3,4+RMIf=C6/g_Wbg-\5>-4Q(-:7X_43L+YFZ&b?DD?M^]PG9L9]]W66>QUE
gEYFZAKDg2Id5GZYc0<:VW#ZWf^Zc<WS.e1<7#(&(7].3_@#&46aI?cFHG.GI_bW
S&PILR>gWBK\1J@6PBJM_abe2R9;[2TC09B-,3+K8(.5G_ce#gZ[,-:bI&RC]?](
.H:@]W]7KRA5fO]A8)R.^N6E6,+X&C93@2<e#6,7c&)P^2W0T/CZc@23XXGZ[ES@
(N:+_L16V<DT)Ag-Z[]AMCJ1HH<DE-OMDY44K(((fe=UB(gOZ=2VG_#QZ80-Z,8#
A>K+g:6DcZSfA?GNUeO=eWLG(2^//fVWRXE6[OTRTP9OP553e,[<[ZAHCC^E64c>
^b;U/IbE:(K<XV-f?4.1\=&<W/,B5aV0A]_F+KS2ecQ1dID.SN8W+/-_9P9Z9?fe
b@F?ZM(KSCf7fV9L?,1f](9IJY1B>/fX_f19U#VN<F:A]53WMTUB?>__>BJC0.+,
?;-J0GB2+VBB+8;Z1VdU]AE@8G66]JB]1gE97(cXAgVd&)EFOa?B==2a?M0WD;^Y
LB@Z6(9FYX2]#eeaBF0N?(dFA,5W\9O9N=M)@:T+7H1e&8-2C24M@OG2\ZNRU()\
F)c4+QH>,S0JFNO-\7TeZIYF#D)<_aE0T(JO,-Pb#M>(e8Q@Q.WHW@@B]#P&1[ND
>YZ0;]?=?\R^>E\+_\L8#)M@6e;EB+[/c/9EXcMX\;YV]XL?><#01R#6d+0T,c=#
Z]#._cGAVfQZ)(:X8#9Gc4KOSGGQPT>_4KcN/T_c5=>RAM]+9JEd^WU#QB?d<JJ4
+@a(G@eE=]cRSQ-=&PeMaAe2M-QDK/9OQ:VIG=2PZ4=0>GDE86M^:D=EXPL@<c)/
+Sf^]FY)W9cfVZ<HeOY]Kd5Y9S9FMe_f0UX9@S/=febSWLA=LP9gEX33K-#7a00C
C<<UOEXcKe4^/aMFf??8AW>&B_[ZA.,(g6OZc_OH1OY3Q0P?&Re;/=EL2\JcXH7,
/J2/FE+5(cWCc11IN8cHL5>2)3cV0+=bPFT]3La^?+#Ng#bX3&P(@e2]4XZa5#9M
NCU7KV7>cS8XDBMCGI-R4:N@,&RZ3B/_<G7aH@JG]fKK58JL+fS+\9J1Zf,U;SN:
6.QHQeK;b(,#]a4&Wa5TTDRK;1BS,=]113(MfTM32M4?(1XGLaLOR_FPc,U5JQPD
=V[Pfb^#64(]ZB/8?cY3FF\7A&-(VfY_5YHd4A13/?(^?R])#E?3>@8:&@SE9f,T
]W:G-?23)-JN-LM5[U3BGb@DQ&J#V8KV/I@/+Cf7LYSGPNTT6N<cU=H_\YGKNdR3
^d(W>L_S(C,CI+]\0^ZP8V\.gCCE]RIOEgAM[/gWJ65f#5\\]QOdNTTHCbE3YcEJ
e7J^?g).H^XVF;<\(M;S?7X<X&F_K\21@UPD?7@+\BKYf+T1F4DDOY^aJDVVSK^c
gXc#SU=Kaa@Z;2F1YD9dK4540?O6@D7\CJ=\MfM3TDe@NZgOS_f<8.WDN,S.BOa]
>RaRPYdRKH69@VLS/M_?<-C8XIW,\cS2D@II,QDa1\IX+9VIG[-CDVJXJ/U2(/e8
U_97+6b8#<@NVV?30E^&1Df>4=eeNefAU:,7-Bb40eUA[UU=127762R5cG3_T&<J
^RKIg@1Z)9+_0QMKTQ7^&,9gN0f<+#SS()?LA;LcGH_8;\_/]]D;\cV44#_K2,7]
.N.B[KP;>N=B#d&;]XS><ae++:f^)GC885)deO.XL]<VeKIaTJQX8--^d20-fESA
#=Q)GWcRDY3#9b[AgJAFe8S^#TL=a8[S>f,27c,1X#/=#]^R^>-FbC-/+-ZS1ALN
dc3cTV?OB#3@EE+27XC</&.P16(\87;NND1]c2A1+;<=]]70Z.d+gAP9d)&861MF
?gG]g&MM86ZPaFcI;ZS51W^>W=bCEB.9[A:(@?6cId2X-f:<?]?6#NF0KF7DXHJJ
_Z#c78J+WT=OgGE5+(D?Y=T)dW@/EB#[;e0SXS3UF@30cSdI@@#LZT6,,PT5+4P8
-ACJN1A>Z<4@fX\-b5a+1^->f#S,dY8W,bXYc&J@N-2,@+6d2Q&65,Y5L1#VWGKg
>JT;+4F0L]eOH/6Y&.?TgKN6.GVN>0K<)F1bBXbdY+)F5H:Z0f(S+-+/F8^Z=##W
@LeP5[Y7)?B-d4.^?#:MNY#;&cY1DgK+.()Ta9E]RR7JU)NP;7JB_+<LYA_-C/3b
VJ1=5EA+WI+?.EI2(@]d-+O]b\^b#KM16XBKZeI.<M9?O8T6a2\ceLO<AeH((82[
+4OO)3E^+T)SVI>cB6U&XRXNX[2PN.GN6\GQYO<<:XH&?8MLZ9Z0b;;<Wc0[<,F<
Gc0eH_/SM8Z)RJb(C)&[/\+&b>:2d2,eRU?ff[X3=3^^Q54H6f=MNM/G?&3Y_I#F
a@]RPM6L<BfY[fD)_;8[5(WLcU1[D+_\+[Ab]ODI=?d@MTc-CH4HZ;N(B3()O_B\
#7NCU&3=^)2&dBVcVU.XW9gEJGR-NV2UU;/IJ=1=WCgYU&P].5.1R+75NYEHQ<<O
,=XH3K<GSKTZ_N@\?I.I@C2;>_a3_SC,AeaKA&JJEM5B)G(4M:D_CF+8ef3;)RM(
+##VQT/6T@##Y^YbUY]^565W3\WUH.Zb?XfYX>T=9Zd>L^I6BADNSH6:QMRU)E5f
EF+9QX@H[<Q<=Lb0-ge@a9C^fRSI&XV6eb0V&GK?^AL(-66>ZfR>5/?\e-1>=dc)
a1+c7\/S:e?R7YS52+@(4F=gObO4LR6]@)O3RWQL5^)@Pc[=^&\KF6:>80+6\2PL
J-Q4G-)#^Y7PQMOMZ6-0bRg]\]99Add5aaM71SM0&7&7V[5_8=LGY;ZC?A3IaDgV
IeG<MffWN)(OLBPA;?@)^LU8Ie-c#@5/I>c+cGU1L86\9A/(R>F7)cU(<AYF51(;
W>B0J:Sb@6QDX.,V,)J66O()ILgLP/ZE=9Q997YUDH,L3Y.2FDgg6E+^LFAHH/;_
]4H1(5.7gTd89\8C11-WXW69gT?-_fM:&@J]+VQ:]>.ACN:OCM>a(()7WgD>.3c0
TLA/+f96+9#f<T^Xg3f,g[<^N.b&,CKeX_cf?MOIMSR@CeQW)]]3NX5fVR?3<6fF
BBeUZOQ42P-K#X-U<@6^/))fW]O.,CE0>0<@,0ff;ZbaU/I2+3c7)>=Z;G(8:S<^
M5G<AB?W^ddJgKFS<ge&]L;?TDA.6089NL4H9SFLYd>&EC,bL]-IX2]M^e8[fU4L
dc2PWFe=_Z219&.e,36bYFLP+4EUD^K@@;D7]0KFga<\Pf5.)-&B_^?F17CIEM4W
2;NLC4RX=6,/^C&A7bFg\[<UW7cF4;OCe,QU3/ad&Kgg1G=#Pf-L@N(\2,+a#HR0
7^QAGdb0NcAF+:_R:5P=SM[GX9^^Z@JUd^c@#FX2f-d::&[Gb^<d4YZ8QJ0^c0I/
:[+ag/CLQF,aM^[02PRP0FCQ)+6U,EG]809VS.B@3YR+G,Z4?a7Q,>/4Q<U:<a[.
0/&K^9+)YOGAHH2Ye&AfH]8CW-[S9K=6gCcf3YM:IBb=;TEM^AVB01J718+cU^AM
2A?&8(@)M.XM:55@F.>/7GGG-gS^&7QbV4]XO5<aD652d:I99&T+/9(<HS1K84bg
,.Y(CMYEb+FTJ:QD4CHT.E8QG<eE?MULg1_eU#;+TB:@_OYW_c&&Tb>X>QVM90>H
d.^PZR2]\>B^gPBfYY=-[@3B6U>SKUT1)LL,0MDUT;NXEOP4?XRCe)<)G&<]dZ+1
&f6CYU&d8(>9-YXKa,<IgYFd74)9D6HP_?9&QMC@/\@1bO5SeKLG<\R7EEI<f.U<
)0T?>g)4@L29e2>c:PaSV,a;fYFUSYcJ08Zc&>ZZR#2D_6?-IYe/3Q3(/gc0?#[(
6<<#QZH)#YGe4@_[6;]g@78/P2fYdP+QS.bW1eGg1fVc&;:Q1.S?PV/gSC47QX1V
6J23<ZS+C/TXL6a;0P85VOT[d6.VOU+H7=UfeY/FPd-3ONU,J3-ER^MaF(6<183<
V-/.NMQ5gN17#@HJ];^<1E?+8ZGO,0AbOACVPTX7P=RWa8SVEV)29L:0a81VgOP4
gRU]&LYG5ZB3N)46(U?&AXJTGa[=1A\PE7/.PaV<c]=Pc+LCbFX5R05Z6)#Tg^\=
Of+:[#dQf@WBV]M&BCKAXTTJ7:RP(0&O?dEHL2=d^Va/O@>&MXe;g62H+NQHd],H
4_<IN9+NX\NR7<F(cBXXLH/;a_RN,9ERQ2KVV#FF=/LdW#&9SI#,2G/6:/J^EcJ/
gA00\ZKK&Db4QB;#QV?3YL[<T]V2K3_]&4=2f0SMZKAV#;Ge/(BBEI_Kb0I(9T^V
;(X(5?Y?0),<^2::DH&W8G45W60=S2?X]H#+dQ&bQOgS3M^<;?1c7?T[^J=G/UaJ
#2B9@C?Z15/RRJ>6Z4L27Yb?,#0a1#@_CfJP(,TS<@-,b.-#8<S/RYR^Wc>]Wd1[
_H.?+ZZ[GI#9\92Y@f+UJ9S=gH-X4+T9;QbV7QR=4HKCCJ4B611\[],3C<8H[c6F
T[9;/:GZAVDb/9IV(US]GM\;U@0GGWC[EP[7E3EgdgZ=3&>-GIJS=D?3OSK\+:S^
LRHK;7=)MGDH/g;:D6@e29OTFDLEJO9HLRHFSAaIB--V]7PeIJ3RdQU.DC.W&7KG
7)\HN&ZFfZRJ,Z=[0f4#C0cYfVb.X8KAS\_3P1-.I_UZe_L(ZNAWP;)#J&ARXDd.
UT_MV1,7)FNN=VIR98@>b4XZ_G+fMde-#SHf/<HCT^Ig83Kg18;;G/>6X>dR;125
K^)RfeYZI+OEM2#=PI=HDQH.)&GWCaV:FL.OK7&U5fcb#18&>7@\M\#Vbg0P:CJ]
(1GZH)_T@^,O<XY/>HGW[(WD6NJ3aTYLgCe7_=P]7?Td-<J?1eSVW)4Q&D>W7d[)
eU3A?[S@BRLI=c_<Wg_-7JHAfN#A:#?.W(eaFQR-aUbO>S\7P)P^L2JCSd<FNKKc
a0g>;;=4\;(CGU6R1?.RH&J06TbB1]>;M(G/KfZTa1PMQafLNPEO#J^YP^O],R#K
C]?^@f2@.D<D3cUW7g0?=\^\9>0_(N_5W<dLHTeQ;&(B+I9,K9-gUZ[C[ZO-\,>9
9@?1I</a09;T7LG-0MP49_fO1b53<UJ(0;-IY[1._fW]I_D8Rc7:<9T]WQfA[U\6
P:NVJCD7aOFS5&@G_+TYdfb>5(H5f4R+d?a(D2XSO+e^dTf;&)N[D.-gRPFQ-DJ0
YUQ#M\_(VV&gJQ30MB<LO(dB?VI+?C@Acg\^<<W8B49V[a7/bW82CD+=5U]9MN)3
1ZZ@]bEJ>FH?E:<WE^#>IQJ\OP,8>SD)VCE,DL1ZA),,=^,c^7a,2OK)YU@_@R,J
:M[0)VdO0TT^B]K<-K:_6_+MfQ08Dg6RY)X[,CN&E4H#XYYC5O?XH@^VOU)8Ta8[
?TM(GXCFPGD+_.BWS8Mb49ge18=6+IY;b^]K2Q>CT[;PQ&0^ODJN@f1<PO\1Mfe=
WLG8[6NW8UV[fJF@JOP>MH\0#LA>BE);URG(;+3MIG=UK6Q=@(\bD(c:8d>1;+bK
aP50\B0R@JObEf&/c:Af9B/+LT[[.RHe4N[1<:_,>\X>UH<8VW)GBb=G5AaI00g@
UG&9eaGQ/>((1E/N^QcAFeL]=;XLN6=@[2DR0(GaBANV]3#A>>?UV?F(;#B)9I6G
B:Z22<2]Zf;[&V&0f7AC4;-LUeEdF(VYB3Y;Jd62aWIF/JS2.Og0I/Gd8W4F8L<8
9U@Z[G,BS5GRT]BCQRVUV=Jb_D1I;8RH^K(T3_-:5Ya#Xg9K&WGNRa@Y5QM\\/b>
D+fE,b>0J<O#8WS6&VV:-I:.=SYHC-:P1K1N@+7/#SBagY1Z:3\K;c3EXN3Y;V6)
;FfZ,\2E6gH1T<J#-.\RV(,dIZa3CS<g/:\GS#_6eL.5d\@>93M+]ALZ[30gREZf
]=/aKLL2LDK_(R<INAP(\@QDd/[H.S<O7EE?)L-7Ig=)/K0[0(+=&#[S=<70cIS]
VbCf=c]7G<1=T<-I,G-/:[H:KgVeP=&Sa:+b;dO^I[.H,#I=[Ge_:W3Q-1IH=dC/
:X^U;T:E4R6DbYSFbW/_33L6[5Z^48^:NW)S#(b.PD[?fLRY\-ZJ_TC?d=/b&-S-
b_M=Df@(G1^3_bV#]=2M<_E)2E5QYAJ^R:ZLS&IH:X(A\.)&,MLS:R7c\fWNf0OI
A/X2FD2:O=;RXF.1),3E4W,LVD>a_N55R?U<<G1OYg,EM5XSWO^ACKC.ARHUa2#4
a5ZAKLBGE\/Z+<aFYPTb8F+faB-6&AC??^D97)X>Q\(=#[S[+@)D]-463YfTg_W[
Ud0(+S;DJZX.N&G>X\/[5QBWR?Ud?KZY0RFPU6GSV(QT>9F&&EA5-P]>HPMEBVV3
7Q[^5@&QX]+NVN+,,+M?1#/c^&+cCR2XO2d&e<AW+NB/Q0.#(Y-NP8f/>0L./WRT
82Z[]]?/)3RE(+54DSK714b3X\X][,3fWWV^cdI1W,+M&JBO_>)c#&)ID7cU<-9X
VT1P0b3;Qfg5/3>DO<dC9WVFH34H9B)QO^DQOA87(&S=IXKUac:734>5VH>Q3ZC/
VVDd40>)C]I+1\fHRbD&7OUeId.0NDf1(3&Ub[E=&]WA,,)Z)=XP5^Z:7-D<:X?;
M#C5UGR[:UQQc7+9e7?R5;7L0J4-_&-@9eA-28.6WF(?S&DfcSBXWR+2<]9=bYec
?4_eA9_PE<ZYEJ?D9,^Ic]#a3YaRg12FfJ+\7YfD,c;RB(>@C+N6F\+60\CR.JYF
\NSD71W[[1VE2.HCLcBTXa<_gT];;-J]-M>aA+e4FNB\\4DEV/4=;V.V_1IR=&17
T07[e>5GY(N+^;\M@UG@-:HH;[;ATF1,f7\9TNI-f,ZNCLR+Y)+[=^BZ.8K_L-R)
XH4G0LY:Uec2gI/WS/-eIV^PCCH]Ve[,eGD.;J^^-34)R#@[^?eNeCT/TKBgB.E/
G&3GI;L3a1O[Tg^RT^Vcd&?I>YU-QZK@MfbRU[IF=E-fdMeFO3UJ7b>5dbT9C5CK
9ACISO17DW7VfA,D\88#SU;\2eRF]gA?HCLNKW?]EFJT8L>eB+[H_NZMb\QTB\AF
9)@BHNC=e.RSG.Y>@8bTCXHRafU0S=UPOS15RCKD7b=#1/W&eQc?TH0.LLWS;S#D
E(/b]8<IVc&211AVZ3RCO;M+T(]3\I6J-aJ,RCS.SU>QE=,>a6d6gRXO4V\/>J56
5=VZ0F&K1G_,X-;7X\cA6QV+5(U[[;@GVTUO@-<^b#&YD2\=a-(@F&8b<<YN,OeW
L_/0OEM9\IJC\GW(:8D]2_2/1Id)Id2?H;^?Y_C7cDa+)PW^>W_RMRg==?fcLgH8
;PPHQg_R2B@K1CT]JLO9ea,.S4CfJ]]=7-JSKW?5^CX/1dNfLD/<4U0<Pcf=.,K1
3WZa+SOELVHWdI=-3_HDW]6H[>Q5Y4E3][1XN>5D(1^\f>=c(VON.X/4<IAf0PX+
bI6H.AC8JNaJf@KZC=EI?],309:5?=3ZV:_U3_2NE3BSR+(<#.d;2HMWf&[R]<@\
B:INMfMR9#-#IWb3&.29M0<#[9F;FU9AJe>#^ME;RS]NL?:_<IW>[EdEUHYSNZ.e
[&=J1CJ^HEge4Kec8[b]LZ3PVW_I/2c:WGL1OQA@(W-G\605\#b)/X)Q01DLGMP^
R)?IeQ/O+T_6L+,RfgIVc,6[fD43A+_RUP<X_IB,K\\QZ[d[^[XQN(2L7Y>PPX<]
_C6D)]6(1LSTFI,a-ge]/b7J]T8(&gcS@b8;O\UQ2RBI5>P+4F)<=>DI]:\PcccA
TbHN+FV^8_?e-[0;HK@2J[2,GCP\?&.ZDV)]I898P83)N6AVNSb,OC.+H>@45J)M
S#:Rf3B3c=9T:K/A4)OCIP,<(cG.O7L-W\#92MFbKNV]M;R^Q5bNcP)d2)DKE68F
:N;SAHF][PSKQ;MI:73AU^aD:;6G3XKU<Q>&^a,/J.HIO/\.fS@S&=(2Y2ESLF58
BUFeP(.2:KE15JVKe/A16]_+-RRBRN>Of4dI+KZT03e1+6U3WHLA7(JLP8+=F=g7
C31_\7K82M>K>fDGLC^>Vd/7:NF0_NR4]JFPcB>b\Ygd-L7I7-#(aQF1R@CTUV-Y
I/\Iee7+&6OSN&<01-DETVBd>F^@\Ef-/fN3&4>UFYQI7\Z0_0IC&B1,;GM,/RGL
(#P7(OQ+X+F4W;EO5KI6_:.C;0^,QPO+IZ&[T1HI_.9bHARgQWV0CV[NgOT<>S-G
0&3ZUQK2RgBCf[GQ2LP-R;#<>729?TZW@RLVS[MLKZcM2)-Oc_/aJg?3B0f5NfG3
4J.;Rc5#[d&GXe#@)+;H6<O3dYP+7[Q[^RQeQL\/K8IP[:TZJe.Q.,2M;eJRa9XH
FV>M^F.:-.7EZb6gI#b#gfGCY_bL[,14(?9OC):_dH,<X-=DcO1=@T@WBN:3S)/#
KU9)HZ/^)XW,af;-8Y.V8=N0e:A2\Md9DF^+Z5<Z#S7/0NRbfb\>4VG1)VD^D.f0
75e9?EAI5;\C>9&I30g<L>Z-R6ePV^5F,Z-2[(\;IZ42^WR3D6\2_g-N=,fD:G#/
.7b,QL_1d:HQ.<V4KYPKKK7S_A/Y\NEL#M]9a-.E-_,U#JRa@)V11,>D[MM+Ta;.
;Sg>08ED5d+fA:5fW.V)/[EGe]H\\BC7bQRdJ+JBg]\c5eGLF.D7+<\g6[_#J(bW
3e[(23HD4P==)1#I[U<7)DW,^ZZcKR:8;S:H_L^,0KfNQ?#.<O3TG<V?.N9<9B1#
3Xe::g@R?PJG-#NNaQB>UP&A<ff4]QX#-9O^^E-+\2X9cI^d(FKJ7MA2C[O(DHba
]\#P-7M<c#/f)H=:KIZ5f2SXINR=HT+?2e571O+>fdQ80C[NT\BZ+DGLMg_0[LG<
2:WH_@71=[AFU@44\6DGQP3>Y8?NFFZ2XL/ZX)O>fI1\_]PB>CXEa(RV\XSF5L/)
]ZLZV@#a4Qe/g@UW:fTg.USggG)/J>+@5=0?2bHBfDG\/\)G@:#VGCe]D](-aB5V
EZ<\Bc>;aONIBP_1YNI/>]1J-3UG;O+.2NMccK84)Z@V[?]5[XD(42.)(TZZWO2Q
>,X2Tfda-d[WM[#-W_7>B6K01B[@]A]]TU17_Kg\BeA9J)XZXZgRWD)D#PdNgY^1
M,JBM-fMO#8+S+>2#d;HN357,2+XMO@PRM[\763Y\LeBDV8\O68.><,D_A7#BSXZ
[:_QeNLQeIXE(\IT5Xd5,QXAd1DcXJdE..Bb4VcC+^LM_b.:L0a=#&;:2SHNDXK5
78+)G:d>G,@B+1/ZSXAO#1B6#e_dBF@T@Z50&2O>ARJID,+D4>Tc\T8XSaF@B2M>
9f&^7F7OTA2[M7SP:_S(XKM0>=UUg?1W0]/\^[TYC/PE0D_I?GW[/e@HFZ3V&KMZ
MQQ[2L/8_GM&+9UbX)bU<M:?TE6c\<:42>IFN:<<;7_AI=c3fN0/HRaA:F<,,Fgb
E?=9:?[?8fO^F/U&@@]467ScA_JWfM.(R?-EaA1:PRYd]7cC@-+\@:YM0ID\2F^4
6/CW@&JQAYUX5-c<b)&YIKObV#<[X5;[<d;77;\3B)8NFDQX_0P1..GG)gUXCW1g
V:+-\^SJ2^Y;R_7_GFbfH9,3-]G]3R@:aBe?g6N^SP:_9Jb<E[,C.>]#+cP;4AZ]
8fOMPP]Y-Q;AV3;GEgARUR>PS1K+DcVc2/Q7.QX-TET5SC^?0=A>G,;A=#GZ>D<6
D?8OdbH3J<W(-G<:>XBZ?OE94P^@&/Ma+38=H25B.@Q-;:DX<]?871dLES(9@26&
@9I=+G-FU0JU#^BJ0P[D-I<>J.9L-XM<QEF3WQ.U3VU;4S13ZSOgJ^=3@A]C)N6V
=((Vf3-JGQdO>@fMg:XZWK3UDG>N;=CA/5#YW2<b&/Ad<>)YV@#<B?1/&A00V?=+
@L1+0U6U,7@a;Z&Z[Y:cW=d.I-V,6c,F\:,aObHfT504IN&Z2Q5^K#I>K+E-?H+3
]3OGNeVXFM6@gVV;AH?fE,1=cAC6\3C[@7Kd\-VXP.>d/e?[.GA:03=U&H#;A6g1
?bN5;-9W<.A-6ZWWa5#-3YGMAA?^S]J5]7WOG7gNfP4.#@PZ6UC3c>3fMN.62.E>
\e&dH/VcGe-3Nc1d(f/+0fLbe#N6B,&.CI?Z=L0(([d:Xa/W(+4V1bS?R]A8N>Xa
O,X(BE6^AMc9e^&/Ba]DbE#NZbgSU#dR3_9ZXO7K/4G+IIM2[g(N^T<3e@OYAc/^
gJ,cW40O)V4aHM0Z\&a7152A.-EYKBUB&4_@3>8]24;2.Q3Zb#]QWEe61(cfe0_a
FJ(WLLW=.3?ZCHefSaW0_)5+PaN-1+ZG.0gO=]D:2#8]V6STA4\aJPEK6JVV;ST]
JL[5277b-;\#ad;BP<_]4@BbHGb+@3U;01UBaPXG)^)4S1]/R<WPKM_7c(#EG=G=
8RTeOJ[#[>7O:YO-\1gb];fHcJ[01O=1JK)-SY#>3K^G2):A[.I\F]gH;/cJ_?MH
4Y4(ETNV?2282S:_>S-ZEe2LegGF(2<O=CLRdZ5:C4d;^\@^U8V.>W/UBJB/&DV&
3?6_,=V^/@6fH]6=AC3W^BgIU.RX10bM6]C^AV_JcHe1S_e->8?F_LLZA.dN^X1.
<MB,V^(IB?#H5JY8M^I3)=c\9Y.RYB^&+dA?T+98eR6QCG96O[d5&2f1[Vg0g\V)
B56Z\X=5AZ,G#:X&]\D.#MS&RB0/DfVLdZLZAAWM0ME)0I^\</M2bJJJP-.F+,YG
0>4b&,<(>FKC9IL)MQ1ITF@R<_S(H5VY2bD5:Z24C>LOVGAWQ3CcNQ)XCADE]AHb
]?,OL2;)C&<Ze]K@7Q/gS)8GJA@f)@D1T9P^2.P#1,=Z.Pd1]H#8[P=R;RWYEaf;
0B6([eQ8L^](/GLEO^D;20,N7]3](\HSL355N9,=K0T9_OZPI-dUYfCbA02P#3:V
;?)=OR/5;2R&QE@QX;TD@1Z2E92[(4_F3U<R9aU@3_DOE.eDZ2eQId:Rf(6fc1\L
gAM,-Z/=0;:N>5&TTZg0]5Z=AUCWc_KW)_UcR8,?AM0P7]=+?#Z9.M]a#Vb6eRNC
g0[Ld]S\Y68^S>AYf8D.(/<BCHTY7-QI@MCgR4QCA?]#,2>/P;X[C?0T?E.6/EaA
8#.X,KW+RB-NG(>[Q8YC:/I5fW^aYTIUS+D42.+BEd+2S7B2c2H=N58:5/\D:[FG
)+gC8(T-:;JSPW?GB9,MLb.E7YgaFdQ1K)>HBBO/6QBO]d#Yc^:9EFRDU[INW)bg
>f2)Y)EGVQ3GDI=bAR/e>A2J=\7.X2CDeSRXF4JQbA6+B;cA<@ED.A_1;Y(V1+\Y
9DWb?,7@GR6P^+3JaMX[60NAPQX3g:+(R@E.^4LI#98RS/-6D4Y14&_g_#W?-LUa
-BJAB1KVQ-A_3ebI:^W7M2F^6A?a+fN>@eFIf6DR).FH<O?0)=3TXUZaPQ+/7R3<
fCO.D0ag_.6#gbR^BM[_VXJB[NbGJ+>97=_F)NW19fg,)T/3B[1WLN9E=UaP[8?3
V>;VFg6#1ETL.,b]XcCZJ_?Uf0L3/6>?LSDPF>?WC<)bgKOSI+LG8A5TZW;eC0da
S7V#H0G;SZS[ON>d:f#BfLIHDXG?0O7/Sf3CE(#\9.cGe@[FC;,>(R6aQZ0gV\W(
GdfP:+YeQWG2[#]FBfI@:@;ZN,-,fD=RSCF^S@@<M5CbI9?4(()ZZf#LRaW_(P_K
DD^6MGK/C4#4\CU5cMa#;UcH_g+bVM;WCbV?VbPM\I/b:AC-\]C6IG043#9bJ.d6
\-/,SYc49Oa:Ge^(H<LC/SfRIeLKFQ9J/CRg0<=\>]/W1SW676\N^(.@d^V(=CY4
_4[?>7D5e+Ad(1-[Lc88]OC8P@4/ZPDE.5T=O5YH9JGHGO=L9W#<=_47AE63aO;^
S7B+Z,\JUB^/4Bb^92OBD>SFaEO@.a4^4SX_&:<F;^+&S;3aQ#[KS9U;6VdCd5gW
.aI@PeA9a1SC)ZGC0XFNXLN5-&R>8+>>S]fUg4BE/U\+JX&_[JN70Xe+deBFP+f0
O;&VG>A/f@-,G04^2D_KVZ^R81M4bCL]UJ\#U@?VV[V(MDV3cGY@V1[&5XBX\EVB
Ug0Ve:cBaOff6E>gX]f6&,]R)bGJ-E]WGMY.3+cS#6L>T41I/H43&(0A[,@,IQ2=
85AO<CSJKQ]N8(A[<dTd?M=(LBI\=0.&QHGg4N60LS2?Tb,FISe2cW(4/=L2D&-.
XTX6c\bga\XAf)#15,+>2aK+7VC[D-R@F+SFNA7^K(T/=_UW>Fd<U[,A,UL5aQS(
3c8=&bbHaGBBKJMRDZJcVWYdU&[UXD7QDe5V/;1;TZLHA^MILUS#=F;N5:11eE:N
I;[bKQ_?8&_b\(d0_30)Ndf_G8fNO<L.0N?+\&71)<:)G+K;24W97K69]=#>W6Cb
ad1,ME9aPU&V23(IMc_.+0=ODD<B[HY/]W_LcJg&M(Z6&0c@Q_O[+1DI1E0>UOF7
^:Wg9/XR[B_P<,eGT;Fg-&PC9;g>,VZ:;e(V41Be+Ud.WfK:8d_c^I2:eI,WI<&G
De0VHdKY->?AF.YRL876=gC(dc:?R?I\94:BfB^X);W6L<EX2Y1dXbN\X(>QAKK8
R1c4^DA?X1]26?GO>RLMLI#.PdK=5/bB.ALUH^e9J5gg7e<W]1dd^f+cI0_#5aSO
<)g8;@,JV9GMMUGIVZZ7&dT&,d+4g<7T;4N]0@dI&_5fd=Fa6d?J4_YfIY.-gSFG
[38>^N0=UI)9Vc,+4#Y)KdPW+2a;KR::@WA2#Y6EgQcKLP6R_RK<)W)9Xgb9SCHP
<d>OM^d.(Ie\AdN,WU:]49:5<F[AL\gCfL1L([cWL0OL\8;C4Z9e&Cd8Y=ZQDe.d
MX9;6<GH=K=;1V5ONIBW>H/f10/L8R3MC=^6O47^NY_AbXgKJad\LT3c;+_bT,8\
\\C#<LHQ\c6_16;&_d85HYU@H^=1H3VK9^-7@M#9a,BP&b:]d8T<\dWK-7S1_Cb3
geSg7^80gT(Z7G0&=^MEDCR:VK@6B4,LU1+EN>)N(ZTJX,G,3[L6ZF5O#Z#Ua30b
[>D2^C/>(2GCB(.QK:WI]TgCHQH,E/76&E1<+O42#J0Y8ILd;F+?XTef??gU7/5Q
3(e78B0\?0&[BW[CFQ/^C,FLIFd^T1T#FUC7A[gZ+R255SWaf6;c^9Yb?0M.AF[^
aE3YA^QVUYHNS)_];WGRBHC(7O+--2]WM#LNTF<K&T]@,.a-]RB4\/0C^_CN5FML
JN[)?H1);>\[.)CJg^e(/L=&DS/9/;XX]D5K/[@,A/A2OALCGMN.CB#4#VF>T[;L
NRS^Q?gUc9JO4;O94JeJGT)a](e/7/K16--K&cO4^R6R4\NPUTFQ-1dW-,8HF3-?
T,L=]P(2E_DP)E\QT)+b;a+CE3,6SM/=\?6AZ>cI,RQ^+?]LdS[+IK]Vef+@<.3M
QO<)7PG69-<Mg8W##J2gO.[>C-GaRNXgHH0^\AUEOZ4eHY(L/UI?W#FFE[Hbb5^5
=T@F;84QC+GR)^P3YH5=W33;\gQ2C8+G;^UMb5eP\ge<faJWNV=TeBb9KRXb1ZDH
-W>]EXKW_<GRZDXWO._4@#VMG.:ASM>R)UNYX#5C[LCOOcRIG;0)3@B)WVbQS<N\
2a);GTA-dK:aN]gYW4J7AOTRf09^OSa=?C]G^b,;3=F^FF6;X>NM&&?HTJI.1L3M
\<4KRQ)KXEK>3cEWdEFSP^&DdDQAeC>Y5]gDSW4J,.Y=#Y/CcS80+-8cMf5:BAWg
3c<@3Y#OA9BEQ5@=@eY(d@W<S\M>aN32C^RMKWK8(,</<a,XgB@R\B3_SgF/T8CU
c=,K\#.-IZSJKD.OE6\>6&ST)N<6fc_.=\Tea:KDVfX;\F5A.1S3R>28Z;BXb9FG
CH@=2NT\:96T0a,?4:YBf_RS8e)&<:ITZ@,4+[O):2O[7<&0I??@8.8-Q=c[FE+]
:E0BDFXZIb1Vd//?:2>BN^LVg-N-0I)>LdQ3RHc-ERZeb&:Lf[bM_)\J5S1O:?QC
c_R1J+QX<c-VK+,/<I5]@&^MZD@M?b;_Le7<X?&Tc/)VFJ,^&/L)9S#Y&9:N\G,V
;dX;IP47&ES(\=Y>))O6V703gL-g^C&JU\(9SZZEBG(C:&XF)FWTUB1KA&[W3AK]
OadY\/^A,:PUJJbU4?:NYg7)Fe)#;Z#DZ\B25dCN9,J-C3U>f&Y\#/M(c_?-M<(<
6-+TAE+JbYN&G@S<Q0EYICL:Sd+T9BI#RB#=0&aY:Q-SQcJ:J.S&C4d0N2)Q=I1<
@&e<&=&DAJ4MM=I.SP#OB?^>5[AYLVNRAM+Qb,F;Rab.5,D?9D.@\3Q+OLZQIWAb
d9<29C:-^@IR+870D_PW.^>/N/e-LSgMRL9@17^,^IRMU^T#bTN/RebOVZRgZ?Z^
d^AUNUTFPdX;U;-AUTY)BMJEB7dOCFX/K.M7[?7b>8WTFL^V;^,@UR7JbRQPAI\G
_:FHgM]79JK)aVQ4bMF+;S/?aX8TB=KC,&=@\[c/W(5_^NPU)B:I?;BUa&,:2@XY
T-CK(Tc8bE;7gJ^Z;PLHVL33ePH0H,78>-]]]gLGFYc,JX[UVed0H[=B90=/(S-g
+HF__4P&<Nc<G2W#;@714C?&S5g;>H0_?D.9:5T-c(F<(c,UT=T;[AK-XFaX^NDc
9EKP1;Q=:I5L&f4F[/)NUAMP&.&>@?TT.g83>d1]USV8:B1.:&5P5&<>60O[9;6E
D;0HJK;SfZJAB6O<9g:)9ALdZH03[CA&WQ=SU0EU2Ea6XR[:D4S(0^H6beb,F:fC
?eB(Q<0@#\M>WXXGSLKYK:BT/cUB\>J[=P8^A,5Oa8V]2[>L<[cY;X5>,O1R@@BY
VLE8Q0Jg,dL:>a=E4:]S8-KTSd?[29?O9&?Y<B>)44(T3HE<c/2]15/?We05RWF6
g9;)<(VN0:HgNEI#b83P>g+AXUdWfOX?:?6-))\_/<W&OI+G/c@@1AbIA+NFB4.I
(dO5;[cZ2;QP,f<9][=@:PP(P^c1F)?dNT^>f;(SdaITc52>1=f&U3A7>]X08d,d
)8ba6/\Bf>RZ;=+@?1<D=7W4,f9,4JVE66:OVIGSf:BJ:@<:_:P1&eD6ZZLVa3QS
B[+V&2TR,QJ5<,RIN;G3eb0<?bR]6--/<7.c@bR<IP^.AUL4M^1R^#Y>>1X[YY&A
:9HAPL^;II\S]PcGK2cKMJ>VX/)4R37Q_6GZG4N&6>?G>.Z^H#dMX:/P4OdW-^+d
DRE9P@>IgP4-L=,WII/T8LcM9e/\\g)]1/7Z5,336OcZKLB<;9H-^V5W/YDW[8U8
Xa9VRXP^<aJ=:,DK3JPFF&5?2>1_:dJF(LG#-gA.U<AL2E5+VXEVC<f<64+9gU:Y
7J3<TK#>TU8[CQ#S2>5]1GBOWB@78FVS6\HD(:+O/^J@PS^PSa0fK_+T)M](N&)G
H@^LZEM?.V;XN1E,X&[N3A\3I1Gbb1@,B-^Qb8W6C3DSfU,N7\,:DS/-\VPEN8e:
GaH,N_#e/@])(S&_RHW0N<)6;52KRU_(.JNR4E7W.+\.Pf0@c;DE9-Dd3UBVK,3N
G:M\][fcG_O1GLO<3;3<0]3]a&^G^)/[Rc@=SMA4g;0598+K>].JD>Z.@U44D>Z?
I@/IYG<4MT6GYe>KXM0CHcV#Ne/UB,fe9<S#c(caaYRf#@A5;Ab,b)5XFE,eg(X<
.GAR6P#V:D0@U=aL20A5Q_XEBIHE#,7Nb#[9\V/U,O-]#Z[CM+.:+054FLU>T-@S
]EQg8(W@<KF(TU.ILQSN0[C##&D?63SH=<1--Q:f>M?eD1]AbZ;=YBfJ4:N0VSS<
9^[V9PILLI)&+FDVX58UFD-SSJ<:/^EC,PX[EA/Wb<QJB\O[W)A>/f=3H<.MBaKb
Y?aB(95TM3V@>TR]DN\_ZRXYIR3[2gM5.FP4[ZKR--dO_IIB[VEJb&?S2@QYBOX4
RL_J&fHDfRDgU;QcTRRD13NU]:@:b?U]_I@Xb^Y,3;5TW/]Q+[D9UOd^+1@DeS9L
D4H:VP1T^,TYC(#KI8X<9fW+QSG(?:V@FDUX;8/?</^F2&OIF&]E\(7_A<?dF/2M
g]LcEb:dX:#(WdOfa9?N_Wc/1ZX[,H^\\]&?R\MPHM3d\.0\2:6:N+[;gBZN7>Z\
91E^9I;L03,YM,#/1NMFaeQ(Q.A.]_,<V1_V@037CWC?BNL1(NI58Z2O37EOP:5b
R7.7[+/C/WHVY&B0]_dUaI:#5&LPQM?/0QLdS9J8>g:.64>Xf1+KBE2LM6?_eST8
A)_,6ZCW?O(2-G)&PM:EJQIBHe^V;d#X1Vg-X9fR(-+?9/Ug?RZQVEfe0;=4@0.L
.R#H?J328,H69V/c^#.aJ&R6V16@T-5RBf5c)PL.^c?[^8F.AIW)UNP.96+?&Z8J
B)E8\A]M<Ia@,<P.-TO8QSMa]a=T<RU=8F>WfR/[&ZW>/WbQ(d560KWR^WeV;(^/
aP8<#SKEA/+DW[GDDS\g>1,:XKcM5Q..G+>HXSN;LUR_LF\D&Z#1HEU--36,,F2c
E+<RY@6Y]H0+=>c0XI^AQ__YAcaBM1CB]2W8bI/RdK,abL]<,L1;L,OXFS<e;603
dMK<2VLD@HY>7?V?O<FLL);58,6)aaQ>CJ<-A8O>fH8HG]>FOCWFMfe##:QK.YD]
XD_S[]3-(HHKI:)_=<28e?4M5L\P8XQX1GGK[+&\FV-c89Ke,f7:V7[)Of\@_eR3
^UbeeK@a9:>GQT;82ggBEU7]\?[YHeW^EIXJ)g75,@Y#E\WZ6f(R5\Y;;\;e3>R6
Q@/9WE>McAbg._B];IeJA@L62WYC^(TfReT?I8(3JWe/a_V^K-UKRAF#+)6E03C9
IeWH)BcQ4>@AE+OgA]ZD9&eN#;e1^/1f1aU;7V]4U]]L4S=bYGIC<WB)eNSZ98G:
9D\X&]JQU>a2UOUJ)[6eIS&?9=FH(8bK>(2CUVGg(b2A)+g[fR:eVN_:;:KW)FP6
UGXD.N<4C#P=[HfddNSX8S7TLb>SL1>g:I6R;>OWf01_UM2d?Q4DADWAWeI6F[/X
gc=d4&]=7aTf9+Z8&0+a3I;G\)[c&=Me#6=#C8866\7;\GL]bMK9e<:M4TQ4Ca_^
Y<b7C?U@fXKZY06/&F-a(+aB44OUT#6^(7<.9b[.4O;+g2#PG]dfDNC6WfXQD.G@
&E#c1K2(6ELKfe[B94CG@]A&e2[;f2.4L_ZT=;g(20[+cV\9.,X7N;BI@0^M1)DD
I4H4f/ZUB5A;LY;O,0N=7K<dSYbR#,NL-5\TIHd(\:,HZHRgBP@^]1G_>T-&,+_.
.-/#[=(2)cB[.(e#H^+<>B8M70c?.V;2#MVF1LLLRH4P[(>&M(-9cD/G68WKN-,f
OPf7:/&QaR07Qe4#cX.VdFN76NKZRKG_X<[Odf;B;UQKDS>aDVUdA+d/D0[7MLd1
VWK]L[@ST0QW0SSAC_6Uf)8XUX^.+]FG9=CJb1I;eVdZ7aZc>2gONbT.gC&MNC)#
IE[?FR\URB@S9/68(<)PJMaD^&>.]=4^XP#_/TeC,<5=RF&\=)f(M84N@JQM60f:
R.=?-ecWO/9.JZ6X>JLa,+_)CILRQAFREXLM4S0A#]F.]Cb6\<S<dM;QVaDZ83<a
a/MNP95<60?A4a&VL35O;JMZOe./;9)0CF[G@IK]K+RA>DDI^5V/C\?YVb.21QC2
4@IE)c;&X)^,\P+O&A2PSfC<gB)FG\:F^CdIa\@UGYMCTY69;G7+H-CKgdG6])##
V:fgA^8[U&b,X]8X@[))VdAHAX9YCIbDAEagJ^e-fKOa]\&/XMR1#,=FF5#g2=9W
NHA3KAAH^UC0?YWfXZX9UL]b/LE@Q24,[\5>@^DfY)XZeW=(QI_A-(cHfJ[[REbf
NCXV6R)7[G&1Rc[5O=X<J8WDA8[4\=G5^,+;55@J5D[e@MSC>,(7I\ZUR-_/C4I3
JMKHb]\]4?<O]cS.8>Ne+RCG4F>&0RcHeCWHaaK0PfZF\9J0&:f4YY.\cVbG?)I<
LVJRM7/=9^e_ZPT)UQPDg-&F0/:8aL?7S-aTX/F-&V@S\3I:&XXeG.U[<Zg/;JY:
:f2MH1/Ra#EBHV9f,TDgS)\(EMJ.78&G<[C1PcD-547a,N3Gf?<;<,.0e8NJfK^a
BIMZfV?SF=)VEE.&,C]]fHJ:DRYF#C@]b0SAJe)N(L[R<Z);_RS/EG-\4]<Z#5/:
d<EW&?\fKf8P7QW/)B<4f1)VfI39.&g5^RO@QCV>+-=M_-M.F,2?ObKcadZ,@IVQ
_,MZ-a(51X6]bF7=VA+<[?&)c+EJ6ZG^Yc9;+PXP7F7-==S#;6M-1.I2=E@PT^b7
]L&Y_ZW9LR328:)Z>==TLTQ/B1eN2B#M]O6cR7+#]FR^3RELUV78U1,VSaB7X@:S
e38+[eFM?<0&V#Oab6+I?N4;d?RZ&M2eB2D1Y69O(]..<XMO^(3)K77\;4aH&9DV
LWdJZ(Q5bJ>8SR>M#S+FMK/JWL(4?XVBDSIE&B,?3S=dS/>.YZJ1F28_/K#4K>/2
0AbE3Qa..>Fg;S=FIedT6U<BPc7]9D.cB_eK;ZeE1)aTS7Ic+T:e,cH9CJeKB>,0
<Ycf?]ga/KC#FEX3dN6?]I(.4#<)(L>ER)?Fb;g_,dR+FTL5C0?NYTQT-;Nf(])a
cA>:;8[<CSX=TA7VA5D.T0JZX5VVS5J=dgTC0)0FG0B0U)PdVL=E?R36()aG/4-G
dGK8)6G_0a(ZOF5e2NJQ\D#<K#8fU/GGeWbB@=Mb[S5:(G9eHZLZ=P>cR#NM@P.C
>6;XIFN/DVF:W(Q=RU8203#OPU]E;->Ic(WBXC8+3/0.W#Pa;cP)&8_QY2G7^HMC
Aa+.Z<,(@S(#19K?\CE,(\,Qg;9VH.BR#UOeNc]Y[GMP8@1+T3IIZ,0&GO,^7ORg
)D2]=V1=2QS]29,M9RLV1:)U1K1Q-(#LPJ&O1.LY<L@F?<J;9(dKC<YKR^C\;)K5
Q_0&c.SR3M<QEe4HUFRDR]T4M7].DQW&8Ee59X\Sb(?V.O/E=V^56AR-\CFP@K4#
V20ZX,MA274UT97:ZRWPHCQZBGGN_WB=E32\11\;Pf)8SeUg(YA\ZL.Y4YecP-^>
R@.GHB6K-?f59)+[#[8@]R9,0]e1/d&M,2WA<P35T]Ga>5E-13e[H[QL\6M&1HMY
JKI5/cg]87?N.Z-a#R;3bH&cP6B9L#1F2YMON\A,PeY?]\c^VKY\E&H6(HVg4+&V
LY^3=()B&XNFfP?g7a,d59RXN<K8CYQT3Z1^SU8RGN;30Y(WB4HOc?])B?OF;b+@
.\&9R]OK]9Tfc\28)bMMAN-05(WXK0;cb==A/>Q96.=YLV=CXI#:ebA41\__PeSM
/E.</S^+;;B&7c>H8JM4ZaP2/=da#Q5.ZRe5(KRF5a/489WDK\W+L>S/dP2e5E@:
[:V_QFRV<dG)AN5F4Mb+>:#Y0Fa_Y+&X<&DB8(6]PNKNM1OgHFAI:G@UP&gU3=ZG
6f[gG\BWUZ)(>EXd_[_ZbN<7IXb)V>3UIP:GB&UDLARFF5D4B\/E_(WO=3Td6O^X
R7Z##21G?[TSB<187bJ30A@d/dMc6Z7HJ8:;&9cDK^T;aT);W(PgQ7^RR#GOE+L_
,:;2<:EfU@PT-Y,V#@@6A9=/8K:b3#eK8N+_[L\_:;^;]?b#3&A9<&-Bc3N)=:7P
#gUUZ9g3RG=+O,Z)DbH=5\M)IR]Veg\a<-DaF9,\-C/PXCS_Q7BG88eJ7>U(J&\a
Y##b8=]c?>.(TUf;9A4aJD_4.?[\3>(O7egD)F#XbST3??#Y^<7:bD-)S&6<SE.B
@WY#_?:;1b\:U7Nb48_\4HOM.G:5<&ffQ#GHFJOVc@HC]>=K,;KXX:7H5[IgLQ2E
-Q?9Q3X4NY5?C#&]Z>O/91O/JQZ(&eY>6)-I/SO^2R@IRaB;EP0QXYHbJX9T8^]O
+7[(4FOF<Y-&H;R+EE-NDcZ><aFLQg\L]bg57R;cP##7?OZO1;G>/A@6(-RN0_SN
E_:Q5-4,V+^/^\^RYHQP]@\Bf<0gO_MRB(77D:@6^T3PCZ_L@E@/>J3=&Z,e>?ab
-,Bf4L&>?/]RV4Gg06F,5TR3e70]cf\dE^[IJ[c8CR5-1a9UYTG_>e0\&IaD<G(M
XD8F5_K[SCMS68^W/PY,+/88_A2KIPZ7JYIZ@,UOS-S5&&g/DG;g(]-&TKM]eE?@
YM_W(A#KD54?>^4\V?O63..XWL=:Q;96?/T;)0VeLDB\?&1_K8HX1BU^=KFYYGOP
[7V.\8dd+-JY,3I34VR17J3I0CPMPF>(/>9P2210;<Q1JBN\Q#GNa\S.(HAb=MW&
C^>f.WRTcK0Xg39SF<:<_[S.G[0Z82TQXV5POO.VQED_&88MA./@6.:]fF0V=eVO
Jae/RLbXH2/Y(BO:WEdEc^A/ZS_@:dRCAU&GPM4=20@\MQNF,^,JIYO54A37C2X8
+,1FfC2c/RcI/L,bTP)Z(^bIS/;/?&Y?_bW,bDR216=geRSK09_eR8/W#M-56F4=
fA72V9=c?ZAg5OXU#P_\YHV])/-@@AbG[-/1N(_]O\L84.RGd^14MN^.YRXRPQbP
VYFb)Q[a_0FVAP1KP4BRX5+TPIIRVKIEP[)QUG-W[QIgF8#g4=S3-7W-K1KGZM0Y
TW9047=#M)DR(-J>TLCdK+Q/H65NUD)0KWL8YIfCYX11g8Qdg3HPAg9_U_/^1V8C
c[-#.,RTeNJ&Lb1T=HKQcC4:f+GBWMUDb#]?1\Te/O\J9J>>]B>:2)1?DIELfb?C
[JQY=ZRge^FH5(I6KOL=Mgc#E5\@8baO+Zg&K7I)N=cQK0[.;+6bc5T_-5cT7FKI
E=K@Q@(O3gMc3FaCY_a[,<\d\5M@Y^6MA,,L><P_;CbS6d+?;R([L4N&eKe56H8P
c4=?8#2G;Fa/I>7@KH.C>BIV7>?@Q^ef+4:/b_F^E7VID\O+Uc3^84gP<>_P:Sb\
DfBELTMOEKgN&<AOO;.:PK1S<:903JU&0O\W[[31aWb9cg<[Kb8E)8),Vf](#JT2
gV3+K.A.O@eHCK2c\,]9O-)UJKcF2Z0A0E[9Dcf[I8&9c[c]PWYXd3CRY&O#c^_9
e[?1L=Z<fIIYN3b_FfG@A]6R[D)G3T.]7a1A8\0Z7S\8R0CJAf\^-QG[<+K?aX_A
#\BQ/RJ#EW/gRU;QK7DHQS>T7.6g/QHHQGM4D4T-3-X_+,Q\e2(6:](15OTMGO_W
,9MZd?>3XTC<NYI03g.7K9GeQYW_&MYGUBc7H@\DILO^@1TT(WF,/;TTWd4=O3<6
SZ1gIQBQe.D2Me+CLZ_M+E>L_T&f\S^YP]0g#[R8H8H0<@BNOUN]4AZ64_#C=F>7
EN1Dg0TVT/N?KH?^aEESHPgH4(5=HeANd5FRY<?SU6:;32H?X&3]6A[I.)^\51^\
<1fUC2Hc?DBaRBW-1B/7IHWH[SYMNT:1\dcS9dR1XUUJX?DK63c+S3dH7W??0KG8
fVP^aS(/REbYc,#UH=-gE-&>8+S_1Q:3(.=R=TFOFd=c.H_&YD78PYLNKH6TP7\W
J1/MAAVdf12(209.KYW#I(KL6<-\Zg0\G#8#U/c67JYGJ&&_+@d\0@CL-L2^IfeM
/6QDFIAH.aZAd_@GP6VBYb&aR4Z?f=a,d=(08HADKbA(2,MYA9Se\;\TUf=12OXL
f>&_aDAVB#RSZVS>-V/LJOCU?TJ)AC=_ODeN9&3WLCR^^cRFX)-dG2e^LU#0A<d1
&PY2[(&,;ZC<+?_RSK0fMbELK8)IBEPRUDgU;>0Q/3[^Z7Q2]&4-Hf^7PCc:WDFN
&/b/9R<.[]RT/A-.[^@9HZ(0M@94c,,MH1L;(1>:.T,HB@:)RQf>Q&#Z34[M->\,
Z-?WXNRTBAF_?XAO/(:.+,#^bPPQa7R^(,)4[,Z0,Y68B\U-=FQ&]4d6#]NZN),b
XDQRW/XT)9XEa3H++WRCQdU&d^0Q>7U(0/;R6KU<;d7NND3eKEGfe,OO#(X9922Y
GcS9SM^e;+aZ@KV4B>^S.W6AR=_+T1Xb^]_Y?/d/E-(4J[MO9a8ZW5GHFVg9&/6F
44Lb9LX_,?b,BSN?Vc4,ad@Qf4+U_f:YNf5?cAb+GP,,Y_e0\53@<N7A7_KQ::1R
c<c;-.BG0&[aX]2Z[S\;#?.KdWSM8,T^.>S>W;;:e=Md4CbV5-[4#Nd@;]8@FOcM
;e@P5X_Id93\C),8AdGITO/4#CbG+LI.X-YRV9Hgfa7PLRB.c:b&NZa0+1A^R#c#
4O82PTaMaBB3)66L-8=@)OWY^B)AXY<7C6EONM/B<,_CRK^?f-Ba?+HURFG/OROD
YV1;;)9Q18d\/@Gb;@.bMBN0DM;XL6>,MN,_9/WN[LKWX^5QC;4PE,Q5f1b;ePVD
[VRW+9:CL6C#>MA4Pgf2CKg^09f\U9\0:+#\^4N0@+3?#cbb0f2.@8/:e]?[2W+)
MR@H>.),L=1-gDNO1.IYL]7bALS;TEbMNN0/B.A7S;fG6PJc5d4@O/,E:da,(>JY
dWe]P)7AZf_X,H,B#TYTAL+ZdF@gX[Ye1Z8-bW+_:(a-JN3+LR3GO2HN@8:VPg8C
(T5@>;cYC&,ZS,+N&d]UF2VV)FISG:E@]XHO7=G=64CJSL25ON9=SB&L];GD]EJM
]<>JO>/2DMg#_cgAQV=MCNVe-LB#R62JHgA23F>P]H-7e/1Dg];L>c-IE/N-0?:f
Z2Q[B\.+=#@EET-Ea48ZT+7^fd2.CUK:W+6B.DXcTU+1K;f6Z.\FAZW+INN(@?S0
GP\Y-@N_ZHZWSZSfCVQ_?&+OHT[-M,=OdSMLFL#>0b\/bKJ]L5Yf=7=7Q3X3bcHD
cTIUTeEM+A)IOP/eEU;K>4:),cF0\_a=CJ?ZB:(F4a_YIS(&,cA+=GS<M:]K^<9:
_C]E/_5+393M_d\7BfbEL>\Y>4N>=V358fW_&d^;cba:Ba5cLe:f@61\+1?MWSAK
05g:0]I+cUAS2XO^[a2(:&5f]WCP<TGY9_8ISa(XRI0Q]D^N(U48\Z&QS&K\+H(4
(eIbKG4K9a5:If^N((7XZ)d_HW:5ZZ<]X4ST]#?4DLB=\./G?8/2(6N0PRNP_PP0
Y#9?d;8WAUPM521(P^XQ(YGR_?ZLA_QIDN+X\c.[L>D+CV:Q5LB:TXWQ4\-6:EO)
UQSQ,>7F,SBZWA3OUb&>ZUb#(ZB@bU+AWU6)DJ#F7YH5H5(?_&PSL4H(b7UO4dLC
((c+7E5Pa&0DRJ>d/If@0IH7V;S-T.#8#L_V33,/F-,F1G82.V[@[_RR?;IM>TLH
WPN#XZbW.f#^H-HWdH5_KR:VNIdY9VZD6IYHI=AO1ccD+BW-RVA6D6XAdQ-0FE;4
0Z+KW1VI;XE1V?P\.BOb6R?\TNPMPB3YW=J,BS.V5.]WX+:gA>^=c=AO/9Y[F0(&
D?-&X1\4XRUPd;b^dB=+9d#/18-=ZfA.V9N/c[9,d7K,E?)P\.3[Z=(.[-Hc^:K+
#UJg_JK30LL0=/FBMF8[R8U8M;d,>IZ?_Z9_NPVGUB#5=b:/LgH]L]7YMGc(^]Q^
+;-?b\LC]Ug^fB:FMFJ#P[M#A4R5>NeLX<.0;G?8.5C)NfV<N5Y?COJ\41TJU3:I
/YF]a\THN7)>Z>dKK7OUED6C;/LF33?CF[QB;S.Pc5^gP^-Y22E3]K5#Eg(<Ff@C
E6-F<3]M>->KQg<7Dda/KON=>9?5bD8IC8eR40-gO)LWC:cDD;G/,Ab<DMR,dL(.
(,Kd,RY[P28\gK688J<TZ8gVV1]/>);5Y-Ja1bA&HG]J=K9_(<:)COCXVO@I6P0U
EMC4P7dIUVB76c3YP3A2<9#KHAY+]S1K@X1#Ta;:Z;)01Z5&Ub<H8?@M\GLD/8)8
gO6e/14RB[+P[:A>DYbV<H6,0F02AdKeLWeP.OAH6fC8ZX9Y]YNc-UcH>a^XWYHU
R1L:JRK/K]e8bB(4PK;#_#/F&3+N14Qbb@&O,YJ]ULVED#eXX\L^#^8R0E_e;XH[
;-U5N37(Y)&G-FJDN:>CES8-eVI->1[W04--2EC,8ZG0?;aZbaX#MYILT1a><P]?
7/].?c2G3M<L38_b0>>D1X3UKR2]7R776FRN;8../7N=E;7OU@+D@CWEN=ePD@d;
RNe7MR,9L_+HHDYI:_Z&3;?N4^dRY\.>4RHY(F5C+e23Q]5ecA@XSTWd_=C[=d#b
&3D25b,4)]N/=ILKWgLUPVI[_HJaIH^J&1-ZbRbG#RW>+&PK=?,Q8d?aJUMLVQaA
XeGB+\WJA/N:9GR:ee3eYD)0&cBXC-]f,A>(4>:&#\5B@4NdSa>e8U8[MR,&eQLM
G^M3LaMIVMRPU-H_\L-Hc5(f&BYCccOL#-Pc\e[aNN>E5X?3UA<39TaI#=PTH>->
R^P[6eCQ=I]S=.>DNJ)SMZR,4b3MB9A2S5.R:BCG4DMV-b60NT\\E5H4[C<Y6d^1
GRg.^Ob:O[.YPH+9c1ZUK+6.GHXS(A[?H_M0>4&-2D+Bfe6.^4R,cbQD-BDC/,F\
,=^P@=-CC(aF^Z_cVRVPLJ?4Ce)SJ+?FQ;4I#E&a_(GKb[L;aSZECc.QSZ>g1;KF
+dJb,^S2DJ.UWZ]72H)DY3CP:/BMZ-&+a.HN0AD@8gU6D#7\L)CBS:4Ga\^1(;XV
##>Ue\YA-LFCLC2U@b2eO^R&0fNI6<\d7eS&S-10<Td3g,=/<@+:]+;8d^YI[I6,
9:86+a^7G:G?2M(FUc^\A\+WJCY-e>QP1--Le/^EP8=/.NfCL7VS5._d^FF\N_<S
:J8FR(O7J8M<Z[F+=:6@Kg5MGA0f=:eQHZ-[Z0-44JQ53Q2_.:;M3S?2,RO@()Z4
b@+I9a+QDI-K82Dg5@&S]W@K82f<TY4:A?W[R2HJ/#O44_AbfX@\<NV49f/cNL[J
;O==Xed9-&WP+^0g3[WAML+F1\CUL-a3+QV5RL]_54W>\SH@ME(KGR+->GeMX6Kf
?gcV^@?78/(ZdO=IH-#KPH?ZKA7206BS[P.[Sg)MDKa_A-P:5:MHK8;=[MGOK1(Q
4@P+V^SF1+4I+N:CgIEYCP(44P8<cbdJ,K6T]PZFR[cdVI]eK==;MR520]&_\+)G
;Q.8RIXf0SPL_7]),.ENf9D.Q^:9^f;>3G3IARJ6M4^K;RaEGL&c&UEL8UKUWD.@
-;6+H-=ddc<IDCOVI[8cPTBN._2#GW]J/]\Na4>c.78?ZU(^.-7:OKc+e)_U2+VA
^=bW3(/d3(&d>24(8D2:V9&YRH/<]#Q#e\@R2)WB5RJ>WTLK@-MEMDeLF_#cDFYI
-=SPcbeCSS6V_M:TIPQ[.bGgYUFg\2,6OR49FRc42-,WYV+\?CLQe[5@ce?T3X3<
RY+PRd?,>G.&@eLJD@A@NYE6AVI-C8WRLJdZU4FX[7(e;dY5+0EAdSPS&?(c(^UO
<V4,.?LT1H]&;gA7P&8?bJA.>[^M11;#LDY@UE9J+\3.D2I?4ESYc2JaYWJI@^+/
eO,NSKdBK=Z/<H^N:BXD:ASWUgE)YUIX2XWW^@CeEJ6\6f61SS2WO>Nd3^-eQP\0
DgKg83K\:?&L9LTGSH9aeG/9eU0F(>_,6NQ-8:#/_U6fTc,(UVH6dX,:,QN;2A^\
M>7YP:ab=I&35;PC,e^X0L5+cIW-:E5W+#a)&:07SD>gW\X[9b@:)REcC5+3eIA8
\LNNORb-6\MR<5W#2-dG-1Sb9\\[_f:K9VZ770T950TK]BWVZfTDE(SR0\FK@GYX
5UGWX)4,:6H>+Bcc>G=TN@<OX2Y#YV-158F?Oad20>?FV0eBdA/NV\PAAX/YFGY1
==27]]:V<Rb@\8RO4RT,9=0]B/f@1eRF[O(XODe@.QHTede^egR9T1C1OXZ/K/H7
7KG1NJe-BUXL+@f&<^A8T8F?D<X:H#\eC,&aM&30^LR;.IL(-?H5BEe+Da.LMRJ:
XXe+]78CY7GGGfKS[.^afe8&(<Bf9Y7.#9JKV5#F;VKIZJ^5HX>ZJ]Q1WBTI=0@V
YM5F/Q_2=MVdEK[HLEF9._[Z7A5@U<JPUGNLMeTHK(b9X+AK9;NLI/Q2B(:NM9^1
F^Y<8(BDgIJ16Q3gV7gb9gF(W)eX-Z5:aaO49<XRcH@#)eS\GK^_9I3@Z587)e?;
&4X9K_Nc1K),PG^e.59K;[0g,AP@Kg4\P>[Jab+/WDeAV5Q#O0e]?J_N>J08RIgE
.Ld]FKUX2)SSP=e7REGKANeDXJ6GKK)5/ebcgJN-5>)XTVA=-<gI8NM[6e2-GO+B
e/[[;4+F;f##K\L6KM:[.BDA6I.N>2TD\D>.2DBK&#]J7=]Q^/ZGa,BV&E4NP.#E
6gae_V]DMN#4Td5U#-?FAW.J<H#2#5_J)f)=+T(G;MNG;E&JBRC1\cfX\Cc_-L;F
8Ja\2Cc?^=[U:WN)b0B2RMQ#V\geO1;=F51X9A28??J@[^D9CJK;C44)0:;HM;93
<0+,Ta;65G\BP4R=@=VUBde;.3NCbMTOXc7NbfQdHJC6W??-gJ/9:@GX&5C,Z/N#
Z-Z#\X7TH,AE(\]&a/(<a3MNB/Z9G[D;RfF&[^L5S\6:;FPE&J1@/?T2A+=f5JRZ
5D&)geX,NE@aP:-9G9?#[NF7+?#eR[<U=V.&4[T)3SP;^44)@6M?#S\<#LIMf>)g
6)Ka@cW6PIM<RTa81WY_HBVf#J5W1S/c#>A<E/dZ]-;PR++F7bS;49<.-M)(V8Z3
3;?UP,Z3:^90ABJH\Xf,SCVB?D?^O^\/V.RY40EN7CUE:(4/7>XIe3C;C]ENE34V
GAYcQ7/<f51:COAH-@aM^e(ATZCe_I\g:P:6E(V>\S(\:6;QZ.LPJ)=_NTdLDO)g
?A<-5^I1-T-6[HM>>[N^SPZ;,#0I8IC1S40SDI4,VdQ=1B7W9DO-]@]0GIQ3#5TG
NC?EBKFD9]4<^bHC8M,PGFDCOU(VE=c+QY5&O.ed1:P64N#J+I0:I68?8RGR2PA3
5.C9BA1B<f6^]_DP;T6O[7DL8JAW]6R&-,CZcQGRCgM1_@?SR3dVU.,K42XHPXGT
M5g>G.K6U:Dg@U,@8+-g7VU9<5[RSWbJ=0&8?G>/XA)^.#<5YI=1BO,LV,TMe<@E
+g=bPZ/F2#:cgI24QW&C6V2GS0LVDM\_[N[RH@#E>)OCW90Q-ZGRBd\Z-cOaH).U
Y4)OLVUg7G1OgV79;XQa5N29EX-,=M6Z>ULZ]7HVPN-J210^MU]@dFf60b_f<=#9
d0SZFcd.[>_]5XJgb[?:gF/_B+d(+1+E=R7deL>Z-21TY&.6Z6QGYaY1HYR?Q;0F
J:(=#ZfTK].Z)HSJ5/T4[VKGD2_Kb9AV-P)X+/NY+g5N+f=,/@]>Y-dTQIF9aeI>
CA>._:<4Pe8\9[#0;e]X6E\HI7H_CP:K6ca-S2Y5b6.[ecKPSMW-JE&\V]a+(&FY
./_Lf.N[=5f;#0_UC^<@VIeW^0:7SdP+)T\6gPR/#b]Gc?9<I&Z?,:,3gYYS44e-
f<fLZ;@NA2JGKSbaD45I3ZT4BEMJO23da2V6E3Qcb?->M_gJD9XAN#V+&V[:K]ba
M?f;MdX8PM3IJ=-a+VZNbd16.,AGA^7Y^?=,Z5Z(5/T+3G\>8^>8/aI8C<G5T#7_
)/a-?D)4OZEPN-G^dX/[MJE\KCUU@gS3L9QT0J>VK\GK2K]?c_8\VaWSFAfU@@9F
fINN33fQ[6\W(WKD3ca>9<[8I-=WBe@Rd-Vg7P:RR5;>TWgcff]OJ4PJ7?7&BJ#4
R-19K-fE_VY+Se)M5+OY9PG]cOWO2W/OB3NVbM9S,eK9TaI[aW>?WdIfZcRS60LQ
N[G6P3&2cG]\T&bU]?a5K&N6GG#_D8T2CC(I(=6,#3b5]FVG@#cb.FCQD68AL#Ed
e=7W\.G#ZCOP_VR(D7N=+C_@A0e/9a&0C4e&=RZ7b\T#L((Eab5a:B_9>2R6)Zc4
:;?-\1W<4U?:\PAD[f4:-0X(BMM&2TG5XXF]E#Y38b^HHA)P2FUN]#4)J[W64[TG
@D/D1O@K36d,ZW=e.2X<^<7T5VV8e#^\HYTL/L.YY/FSEV.O:fN4CWR.7#,K+TJX
IQ?=CA<R?7@(=M]ag6c@.IX&.1CM(K^S:05Cf_T.#<7Cf2W=&T-<,R/PYEgO49Od
,A922:9?G0Z#da3bZL;0OSZDDcCD&AMR3<aJ-JgBUEKPJ3^4:<56W+AbP0AI]>][
dS&XU#@,T_(f1M[;PA4QWQ?3.9gRe(c6TXHW_7ae^CLT;d=MbR4WZ&Z&O#I;#XL:
F>44;CbbM[F1]^=VET=JDG_&H+#eSPd0&[BE]^<XNMS#&e[Ga6?]>AZHQJLHC7KZ
XQUA_KQT5,/eW=>W)7C_^0UC)794,bWPI=8U[\,26ND]-f<.B6;+cGJM+fg>4OY5
6Nd9c---Y=Z@5S<WB,NST<7+)+,db64FYTWZ<DfWM<7?V\IQaN&^U-e+?.NHJ&.b
Z&aH,_:FD#cfBX/6;d_Aeg^5aO2W<I0H5QO5^0?@<d)Wb=<9+ZKS&BDb4[Z7ZD&c
dgb@Y/,SfG\-BP<Vd?Kg;]eP13P.D<BF9P<d7V>.281)9[@e=:5:7a49efUe,M^g
)48WPJRX]FQ9S64)3H>)H0-CV^)GY67UYWdYLUK6F9O;_NZHS[?&cVF30FGgH?Y[
c.QQA9AM:NgbZ2SdWF6-GRW[a#8dGXOKYJS+T.-:IXbIRBGdWEI?1NfbJcX8BQTX
U@:ZL0STU?d1Bgf:VfI&XYL3]MJKSNW\027AQ9(g>H4TD13QQ4[#?;e?E[bN.R+4
<45N7L0H@<3DCMbQ5PSG?1G?H#TE4\ENKb]=@?:8CAWM7SG&,Y227e[aG(;^1ggf
-Z?(>VS-f_ED.5FM.X-dW#P--VQU,@a]cFc6NP=&<WN<(C^ce^<&9eOR6NFNf5fA
cQTbKMfK0LLQ&EAVA@F0b7X]CQ=5I_Qeb\3C//&F&)E+(GQJbLI8:7E7#4L0U2ae
\6QZMWP46eC<7M2A?EccccB-AZ:a(LQVF,RXIF\W,TbG30S<WW/aQ,UT)_MFJd&-
:I&J1A]H+9#eH4]/81KBb7>CFQa3)4AC<3&L;^W5Ze5#J-W?a7HB6R+7DgUWObO6
8e=AZ^1)3(I)H7(H>PIg7Ea+^\Z@1=;4DI<;^D;IK3#Vg_LK;eEE.DG7V1BS>&fA
+K:?^QY62C<_O]/be.?fNQ+(TQGKM[RMD]1#3J#MQ2^&,F88VFN/DB2HD5ePZ689
NLFWN7@)?5T,MdEN)_(@\2N>M:P9^8@HEa#1b6bH@JA3I[]PeL\9#\S8Q-\/5]7[
6Ab0KY/^GeQ<?8O-5:K<)54eXH&8Xd]Y:NcD^L8a^20FFG:R+7IT\=.AX6:RK6GR
Rg6/V4+3-@#H)6MDNb1Z)UC>eXI(V5/,SEf]I,99(9b7QecQOL(8&=\D928QMO+d
:bF+GS\1e#1^2G8UWC6&,Y[WP<_E3R0_HWB].IW30+GL=SXO[]EGJNU(a(>d9RJG
1fQed]OU50HG&Dg^_]5.[R5A\F,:H1-fS2g<W7H4+7A^4>b\K\9ZT9C?>We)1RR;
>EFefL5P@^30Ogc#7\79?&L>fKF_SN2)CY-O9g8bTc>O-5ZD9ZP[/@\FQaL81\7M
=\=LN<\U0=+HeT(0a<2;4/<d.e0PV?>PV1Z(QH3BG+2fS_J\gH.G]@5QWO]F[(>P
MA&7I9D?Y(MY&:U@Ja:-dGBGGdD+A<ES<RSbV/;TQV?E\@)F[Q2^FJ=LF4c;4=+I
ePM9HWWZ_0ESWW&>.EEWF3H4eZ-CV\^Z+g>U1GE/df)QU,_gb=ZD5<<E<CMc+5gE
[MS)@d98W.839P8_)Qg>\_d-G.X,c\LJSU;YA_FA^1J[V,-ILE?C^Jc.D/e16AHT
5L57-5e78R@1[13TF<gCA0>X+0[M/_IQNE,d,^E5C(fO<g[@5=[N=Dg]4&4)eGI8
W1/95\F:VOIA=SC42dc.Y^VbJgX43D^UDR9Jg9CV-8<7dU[4R3.+WCe>]=^c_DJE
B:8gG77XM&RY;\296-g7L7/5]0UCQaeX74?eM;L]QA11-CFBYCc[N0XS&3#?C\c.
9eeN;E)Te.R\E]@R6Ke^N=\f<3L4S:M,NeIC,F;a?2ZB7Y4.33<07eY/e?)d:].:
.g[7XL(\31:5.QVCNP/0L34LD^?GFNQd7Z<T&5K=^g-2([:dF_T/OL>>f_KQbC-.
GWW-,3P-a[@/I,g[.7FP/RG;Re0FREPJ&&/^][0dQba4S7Tce-<7+ZHB3L_[(TdB
?a](0DZaNgO]-3@2+GUJ-GUIMZcS<FFDA2,4U@1JHW6QX\^fe<,O8<ZLVXK6-L,5
d;B0ZTV\b;<MS)P&e+B2BgYc5?0HE\XDgIL7&&3Tb(K&[Q][dKECH<RK#R54^eSV
fT85P0R-Z3KKT@O<;V>AH]PXUe2d>A)ROgRe/;P11[&_2LCYY+U,I)e8V7G1JQ#9
g<6.&,eZS5P<^4NZ-M,DN&bc20Ud-Lg-50+f^E8b,8OV[(+H3W.?QHJ1O>=2<[&f
_E]I@dF8Yb[U.;]>7I]J5b_G,6-J84a3V>A\;d:)3&Aec\2O=^8[;IUBB@3+Q\MY
+HQH,N4)&81fg_U@15=9\1(XI<W:B&FOV-O+\>X)9fP9GNc62^XA:W+<G#O=_OK^
]b)eNDEI.Gf.a#<deBQ^)M.T83\g[];8WQc]ZD^_:XHa\NPTIP;7,X5R>0V?BSJ)
Y]=Ef2]7c\W-?Jg0G5J;fLY300gWgCSV\AV<dNYee.><H_^?3?F2<S#g]#6B@NRI
^e\4[;L804Q/<P]-A?E6d0b;&3bOHfY=.]\BO?S<a-b19:baY>>5E.aE7IaL\af;
[QB?RA1=Q[?9+]ZQ@FM(P-UAP8ZO=Pfa[Pf3^b3NTCGT.&?BNR-8.]>2fEXI,.0b
.ca,/^@>e:/F6OYRXDNVe\6L.O6L=C0+4J^DF^+gR^1c_FTK<5fZ;_aV]8O@9G3,
aAT<5-c]#S#O9+B=7FI36Y;\5^&A\e5S_BK7&E<eAFc+G>?cJf,[0>H-EA>;PWXC
X4?e2NULZ)FLTcR2RW,@=B(M#UD>fb0P^M=BT>8a>A60+L7a9KOgKUZ_/1OB&47/
8=S3cG607GccE08DVQW2^.;5=FG9Z7/D^8[SRGH&=F:PL5aLY6V..B25)McR,8@K
,I2^AEBN:N<Fa>Z#SfE<Y=(Kg2G0O\bT^NF--W,;O1.[=5ZSe7fF\W14aKF_>8[Z
)=;789c3QUGRHT84ZOHRUe]LNNb5=]T6Ne>PRcNE/E6g#?QROS=Z^X^9a)_>;aY?
;ODBdH<3PF1/:R[UU;DXSPNMCb-:M/]f3/?Gb(1=-a[=>-(.=J2X,MBUbK7MfR++
(7Yb:fA.USN5FPY^0D.S//B9=0/K.P0/,Q1XH7Yca,G?Q\e(6RP(<>D\e+DVS/7[
VgOgLCS]b(.@4TF>2S+3E.L.WH5dWXVSN[:aDNWUJ^N(1QaN=#b0E[ZBWQ#Y5K8G
C//57@VO2(a.IJ.-N+\URfg&^bL-8)J3L[_IZ;V72bfK>E7V9.W@[cV,:(_e;cNR
BbY]I+[=BGW,/^T39Z8[9.D>eWJ7LQC(Ee&K?dG=(.2fG9&FY1;#;=d9M^-g.WRO
)4c723BNBfWd@d4gQbS_3GJ(N@P@ecFNbdBN2J63?.VFf3._gD&01W)-^&WB_4C:
<T3[@dLa1+Z>7^caU/_Zd/e(KW-dZ0=X_fF;?eDI.\)V49123T\Q3#T,,BN<=BV3
3fCHgU&CEHH[)BL4FKJ2^@R4PUK06Lg\>?DQbV^&I._#(3IT_]NcV6=^IWY\VSag
;?>]EccN9c/ReUHC<^g9#W)^7]WaZGXf)6a[F/Wc5_6^TMK)1gS1(bF9EEW]0EL:
P,L;g5)Tb41?F58,CRRADV\Oc/.C1@+0Z-3>\[KHJ;:eN1]35<+C5;-gJMa;e(Xb
BH]VM)a&25V?AUHQ:(=EO][V63</gR\9b5?L1P2A>(LWJO/W;].KH&DG;WC&2@W[
)Q0NVW=P\f#IeB:1.PW?7M2X]dBePXP.I9,fV#R85EA0)F.VB<1\+.#YKaX9daF1
<#d;9:MXFXDN9g91@:>Obc=C0\H=^U-]fG?f8.PT=4G)&=O)7E?G[S).?^ddX+#5
KY4.dG;.9VXQc&MeRE@;WMD7LeP+PgUZU(SPUFERPA4b[BQY9?:BYP<>7QYDgHTV
d;7ZYT]T>f\d9b;Zg:?eWC?B5Q^:PRdgf3S+<2L8Q+LTAf,,J@(8Q\_0W.67Q(QK
M>/HJJ4VaR^04[Y-bffgJ4(V-_#=gIN@Oc).cTNADLYTLa)#<@5=TfV+[&47]/VE
#7gTD^SCe),B.1H,3c;:]7PbVO<;54Y;]&QQ3_+^/5)2U5J<a91<2SWdZ1[^.4K:
@X_@AcLD(TG;QU\TFKY?\;TES_?\aQ=YDTdg.PLZ4e/@^A9/8RDVePYMDEQ+;U-e
0@e2=,QeZ@@dbTTTR92RaAC>J+D[A1SC0[VM#^(2<1\.2A\bQ3f-:^\/0A].^:5d
\12,?JAWZKPVMXfCQ#.2#N2ag,\AbLH:GcH_0_/\a/M_cX=WR/==_d?,]a#B6)dc
@OcAK-6)^?USH7>C1N8f.;O^X=H#)U-Ve+2GZLf>[(^)92Ad]H-gRH44@<PG&eDc
WfbQDOTL.JR:O^?>KX0F=E25VA0aY[,_-_+8]3\IX26&KG#_H2>TVbPFXGQ:7R49
@e8PeR+.\,3,62KZ\)>/bZI\B1[)0U+[2?^W1SVPGDdF?A583F61,C?2P1f@?V\.
2[3eIIZ3D:aY<1gVS?NI<,3]Q)ZHTI\K>]8AB)3EX+=JG6Q<LU\@2B5BDUS7)eGP
1G]@X(##RSHfB2[2,:<67ZH_cI=S_FJAS6AEcS,Y713.N</Q5FMSHV0P9.-^RKH3
H(2UAS_XWM]^d54-gb.BfE7+PXc#A#]N>/Za]/86\?[Q]I.C.&>:F\5\KLW,OCdL
NTXQMX.&X.cM4?W+)V6@-F))/.37L#[b9Fg#BgfJfA?TTQ5@?+fRRH^8e&-C6Cf[
#8XeT?R_;M3#(?FC?(N8&Ce;)2XbMV70^MZ_(aXc@dXCL:0[GdYA-?X38HFBTb_S
4RTDZI1UKUKd9OKMaCUG]Zf],cOc^Vg--;A2Y.QZPF-T?>FaT>:.K7W6DH6P]+\)
bE47)DHgf&4gU;OE168L:063XQG[3;e+Z61XP1/d]WXe&G1Y0O0Fc?<HG>IaF(?+
1.2\5@gMEfDQQIYB[SZ;g_3eSQ_NPM?#KdOeW-Da[_,XaFH]N_dART2C+C23^?V_
/BK_6@@)[^Q,@Q3O?f+G\IX_G[aE21==&P+ZeJ@cTHX+fEe=L2dGC4PZBYY<14SL
)^QN14QNPD\VMDG;d8d4G#0Yg8eYQI_0;O0<XX?)Bcf)G>U^\)EZEV8)>T^g0H1K
]g>9D3P#Ne\_4fO8=[V\K^M[?B0/=QFI;HK,#98S8^M\-N(SLRRH61d&HQJIeNB,
QDN+PC#V?HHeYB]b5RO9,#52e.>/Q\S3.)bL_R#N-Z+4\2=<QPQ&C64YaXUSH+T]
(R216d8(gVM>+BLIEgWfAD->&^D35GdMa6P&,3A8QLM(18De_<Ggcd&&2<-M2H)#
3RUH+^bVCQ2=9_W_1b;#U&@X;-B#fR31Y-bNfUJB[O&-1ZG7YL@9B^FT5RMG[QZW
>)eGc0fG=g<N0SO6F&O1QXTB5=V/>>Y_Mg_e8MVH5H>0EX@^2bM8a5(f[aQV5EL+
JAKDU5?E(=;e2]?HQ=6PdHdLK_DS.P[8)=HS1HcZ^NUf6OU<5TUaUdb0(9_Pb31P
F>@.8.BG@92#:6U2+:DGI/87MZ7V&UUd=-UQc=61R<Q>L1UA5DP\EDc_&4gHZI@d
b_Q@UJT1C;(W7X^?UGC@R_4>41CGXQY>^YHETW2U?IC,LXB963?QB68^@G,5S;:@
IRfbAE;@XQeR2^V_<TNBG<G_T1Y3S&G=+9G7c>?1gSG)8C</HIe/b6SEC;<UCNG:
^5Z<E1^E#SHV899<L3Df66GH+OcL>MQ?+CAHTSB@JNXdb6B3[PE\(b<N>fD:G.Lg
S@014.[-[.DJ/E8FBEb6#D]ZgAfbVTaN&S&S]Cfgf3FFP8+XF7[NEXdF3PH@UIG,
E)c><bIFbQFGT>^e/>]M&MZ:cS9dc]D3_b=RWbN95UfSP_e+CgDA49@L:?9X>c47
_Je^B6=JZ^2#=eg3DX(_^+S4FX^S;Q)C>1U&[Fd1^.=KYV8LFAf8aB?NaWe>fcO[
.EAK<21&8@EWe@6OL8RR9AI6J0GP_8]C]8dX2K5XC@ZC8H8gHa#Y<^He69,TQ4/_
S>aV<OD+B8b-_2Y-I-JD282EgB;S)OXg+\;UNN)#=?G+?]/N#/\DA?E)UI6DSJX0
215^-UJ&WT-)4<2fVUZ=cXUfVI>)RACgSQ>g;6dBFM;6FRR7N]4b0GFL34[:,+=1
SYB9W05KeB5fZ>W0[?9VYI90f>C#e)NKV\7/6RW;@ab/80YETeTa0cHBe0.ZfL-Y
M-E_^2U0?.30-73R6E)&RY@(JDW\0C2PZ?gK319f(F@9GELFeV#L;@8LRNgb8H,-
gK;ZI4;YWBK0)QQQb6,7G1I.fGW&Cf[QS,]EY6f=\c@6a=_Q&K-B(a-\LAF?VSD3
TZeBDS#Z&]PA@>+[MD_<0@-c?b9DR0.[ADV]?:Q1X.H#_W@O1G=UGa5W,&9/J0IY
Ya9#C]8P5NV5J[I/H8f=US>b.f,+D+@:+^8?V=3bTb]U9#IcA]&cgQHWdWc.V^?;
fCg\L^43UAE7C:6dOUUH.g\<4ND],M6NG9.BAdd(H0C?@1fRQ2[NXMZ1dC7dH#:Y
QN?V<^0:U28[]gW::b0]1FDFBE,VYOZF6H<+cU/dGN.,Da4>=2VHJ[Gf=\\Zeg&(
c3(Y(X)[]HaJg]O0CW(XN/1f9Q\/^0>?(OUYS>7bBRZBTCT1JH2PMOK)N=GUdcKN
V.dS.f0?.b>8NMaMd]UV&MK)TN]<&#F]0K,_Q79F/>Q@7U1Q5FZ<F,ZGT>+QZI)@
7<GX\YG=8cC^:Td(Y.S+e9=8JD[6MPZE89g989LE>/]-DRNg6cE&EcT(FHT\:\<H
./)C4Y4]?LOED[I)d[E[Q#_LAB=2DFe:_7]U\XdK:CT3KS?dK3..;@+F_RUA5^-R
X&Wf76b)P>:bP+Zdd2:8-LZC]@7[TA2J/OGR9IW@Zd[Z1Td1VFA-Q8b2dW.BCA^V
[TI@J26dACM))?JaSRB<VUY-.)3MfMG[M[>Fg<7VGE;,,0@832JZ+\)>053@4B2J
;ae8a8TMKT4+;9OQ^;]CABN2,W4G@d2[d^7ZKV5K,;EE^^Z6_=98Zd@=QbY3UX[&
E[#^-E)AaO1a&1+-:HEcIW4MBG7RP/g_/,c?>)MZ9QO(M3a64CEaI/:XKFIW;b@7
)K[?Te.bF3E-H@D6_Q2+;IW#HH+OHf<B2LMFESDZMV+8KNI\(11,K+K+H-^]eMNM
6AK;gf9HFb>OLM#bS)7\JE;+5>E6B/LCI\/ZIdOIRSBB^5[Kc)&0^BWH07R6CEV#
EI=O>O;O<6O.)YGLH(NQ?eB+I+.(6,D_dL?&U\>;II[7QV=OX4c@P\UVIcG(U[\0
c7Q6e,OI:U2WY</48_^#(&A\UYL8I@\FY=L1;CAYa_[:b4<S9dcX3W0Fe4?2B9B2
<8R;(=SeV_I8J.3@P7gFeM>Dg;S\6H^L=Bcg^.g?I5+/VXGITb-Cg,?7Og-bGSD@
+,E9d9D8aR+]#B4ga,7J;KQ:H+CZDXb:96gH)5E\6^\A2ZUKP\6Va2X[M@-CW@g/
aMP3K<:H.@fLJdA+PCZ9,F,\4@>)FC1&8;<38gD>5)dK6NafZbS22S^TZd<KJBF9
8_CZN._7W4>Q)IVI3.;E=5;+7.^OAeGG>V]=Jb==9\RcFSN#+1cK[&:VL3\7[Ead
ZgPJH(5YM6CWbg)J9Of-,=_6eS\S?JHT/0J,b5O/edJSU(cJ)W.=4SgB(V>5NAR\
5J]\HeA57JORSLI_-4=H4(:AK<b>?[&aC:SM/9H@FM.fW,>C(\O?G^f+C<@>F3?c
1XM51^L.JR4d2+e<aGg40C8EK9+#IGd7;/HPY1I<=f9U4J7Q/2Lb,TdY26KaK8aQ
Q:^-<]Ne<=B&YOGE7+ca9-;aC\eYY]0HOXKHZfQ\M).bd-N&U_R=K9c:OAYH<2^W
:3c^cL_IFQ/#T2A0SZI+#]46:YK@Uc>4#._0a1VC;b)9d;@;V2?4cPYGBFHHa=Vd
(RgQG,80&51QZGCL;0=U\e(Y<<R54Cb_[_dD\_d#3ZPd9=B&T]LG1F?-NP@d>5bg
0V+d_WJXCCAD/^8&e36PO_#dUF1#?J15,O@+2E+VOUYAe0PKaeQ]3]3S(EQ;CR+X
XLG7JM7VOAF:Q+Cf5,WR&AE@]_Y/RMIKNOd5>1RHRgC+2c6)MAF0?@eBH[2Gg/.R
]Z,3XbOI_g7M0-#FGXTH+<J=#6OIbJT@I3BeLEP1#BQ;;[d>WfS8B5072FS,=RW,
.aRQ]SbMbeY9,+D/#fB0)4T;@Ze;<Sf1=RIY90;#9TZL;L//80[+6=AcBEGL8Q]N
7/P-OTcf]KAT5fLRGVLZdgDK6ZEDU)-abeI65@H\4@IS5R^+L]PK6Y[B943_8W_Q
SHPc_OHEI3/HBXRG)+F:5QYY&.C]Y[-^>O>f(,bBZ.5g)3GH^M?Vc&](YD_SVP0>
BeV<,LPHf4^EM>LZU&@@/2Re7.e1Z?6-Td>aKD+B\+:EAJ>cQ4\C5D\RWgK+EcN:
UBB/HDEY=dDbQJ>U21c4=H2KcD_2SJQ^BaE]3]TUQ#_b7MU;Q]=D1:[CI,F^Bg@W
;fWS]-<-)O21&M[H6@J/6U471e5UZH_)D2JALS?NN>=<FgQ-^IZPNS-7+A_4[ON7
2#@N[#1/eW8QD^NFN0<K>B1g]b5S)J]B.OEJU55H.2.[Z;&Z3T\.B27F?VP;.[C:
8O9H_HG>g<CAS1/0X<A_ZfCX@U.0WE/(V<b(YH)P1LeOC6V&BM5P?\0_8Da./.;L
IadM\<M>LB6.[W^L5@e+)K->U4a[e\4bGUJ^S;2/7J..QVM8:VL-]H2Za8+RcIZ,
NTg/](4O]f<b80.BbF_G]XJ?_TZ,-/31AJUKN^@0,9+;G]I1R[geD?=\D3NKIWgN
a_@8::Ff2WZF(Z1PdCM3^9O>bL0Z7]DFUGK[9EY]-001/4O7LQ4G#XI\eK>)C0P@
79^^WU,JQ=JWHE,.fO+9WRX>-7LEPc0b713E#c3#L(Z95_@QYCU]>c/Lf>/+V#5<
cfMS8,2_ca/M_<+AL,)\(8&OA^WW\GVP:UFSFfN5Z?,S27JV0\CHV6]C27;7Q1#3
aX4ZHK8.1_X)H1?>.R<f/4552:Bg<P4@H>RY#MGdBJgC:3TO0/]+e4-W]a(]7IB7
?7+P\(+Q&fDJNLLGKQO9F=OKPJ.(A1RDFMXdKbK-(6[4(8#<eI1O;X;>VC[[TH-K
]&M]CIG\.40#XP8)9-S@VEJGY4XTB(V03.5cGWM;QN5f0AHX]1EGSff?L6P2_(AZ
ab244;JXQdQa3<7/Q,0.PZMKQ=fWg5/S[<YESMdR3^OA6aBDaa9Wa]V]_S201V36
5>dCOVZ>g[39eY8OWXG8HcG2AY?NE6#bW9TdS;PF3@Tge/Cb-_>_0DB>HRV_RE:N
MA2L,&PQ\cDHfD?)a2CEW2Y&(&C_X&d648[ZB@Z@)^2+)?=d9063PS:+<dAEgGHM
LbT0bF[KYJ7?,@0H(c.>@/64X/A&QDdA7?7Rb>/><O?&V^4Zg2R&8Y1C952RJD3D
U&9Q4:\WV(WFF]/\N[>9E2DI:D2V,aQ55T()7Wd64;cf^W1P1a:2Ie&C)7]9W@=+
I9:4YgfZ]/A^\KUaH93BASXc0W<Jd](UcR&-ZFX[X&KLT12B3?J5eS[>P_(11]47
G)(\aUDUS@fVOgTQUDW:^VZg_,UHcecC[:+0_#3WZ>_I_eXO@J\H[^M9M+;G5?bC
/B\<OZ](VLL\ZTEQ+ObA-.]<MaZX]OM+26.c(I1_YTWE0E#RE0L3BBLURP2SN/O8
/ObVdES3RDX89UcNX\6:a2=>dN2M)AdNcfd>8KHZdLL,ZE@dBXb<Ve.9X,=\1V8C
]g3<40-39TK\cL6VX^)I8]#BaXbHdAD.<D87US6@@?0dHeZH)DT+FaBfKI(0Na=a
Aa;>M):a,\)ac:/2\eKa<XI&dWW42cOQGL/_,PM^adXdf(Q8Q3M=eUBH,(/FR84c
5bQA./&_4R\&J;dLSJ4\H.^5d\>P_Q.7;;.AUBaW?d;;f&=.:KR)8/(4-IXTI3+>
7B/>d,2>K4-2b@&PUY&5^XX:4JUIHT)(]WJfc5f=4c4eJX>C)+=PI(X-9Y?MVWfO
CN70bVMP1IK3U-<<4?-bX5&VG.GQ>8Qb1S+RcFdeKR+(.U6YSB18>=K_b4T#Z1PF
5agU)Rc=4#B-LEXZJ,.e9=.M=#6?47a:gF[+R5a=I9Q4[MfG^8_6:T+#DN4/g@C,
]LJ/WKcHeT=5FcWG>XKK]17<9;(3]?5Fd_-6-I7[@fZ+^,ae.Y=U&__b>?JQc4J4
e<<NdDVM2^a4)D,P@[Q-C?+>X=c@<O23YS8:Y#VY<7IYIS?Z[L:Oa-1^.87_OPW3
>;@[510AN&T--9L,<cT[)(R,/b<9dSQ(-RW\22MF@S>4d)RV-BPD_CV)-XFFN<TZ
+NBO;6;>;W;.=7@PEZT&?g,TG#]H0QIHE6,(bD?VBOJ#5NFN\e,/)EZc47bCZ#Na
>M:ee@0S(>\4W^+OO(4WXX\6E1<5DYR&Wg+aJ<#g=8)4\,,gTZ9?BXKBI8P5A+O#
GEY,H<?81U_VZRcFD:&R,&#VNaY+L0#-bXS5\f([L^1KK^+VaD@GVQK1UJ29&deC
RbU]>)?-\=Ade&P(AfB0Q+4HEdA=@PBM;=^#HXGM(X85W-cD[0&^JU_Q?1Jc<:V#
1Hd0K08CFNF>+d8KD4H9=KMeJa^I;+-DKFJO8BeDI\/31M6-<G6AW#@NYLb2\.6[
N3@2/[BNMeM5CH/JQe0fQ6@dZ-J\6UgE.M<a52\7B8;N>\SDg]QQ1EVHNJ:+.6W3
&4Vf=d]4DIXKg34ANV[5W8WYGGUHLLU\HFC0Qa6.ag5eMQ;Gg^=HJ\@A6UICVgfR
62@GGbW&>TD9eba7#6+YVg-/U]255T148:PQ?YFUK,Z?D5>ZT2,[@g_#&V9_,6TN
[Na__a@TAED^H3+J44U>R.^HTGH@@2=)gJ?)c,Od4[@Y0?IX@6\CRIKIU<NPH^Y^
L6<He>3]ZEYO[)fLQ;YJHg:\QRORK6C;VP8BdEe\6>4.bJ3/bgX\T?V^.-M?&Wa1
Z/bN5Z7gN;KDJ)=@Z7->W\)F.6.0<P<#URB]QHgVe_@_ac[JQQ1fYf=Hf?\)]J2O
SEG,18NO8337^6N79g22^AaH:84/29X71W_5=f##;9.V6485JYSN@<I_EQ9MX@GU
Sa#AEX(6G<fZQ\4[^ZF#6JV@NMagQTJ=EdB\2W]bWD1C&#&WKAN;+?D9L(U-+9N0
E4eFIV5FX:Y;\1.FB4[@<=OJWY\39TND[7M[E<@?6@C?Q_bC;XLC+,X3fg]T#>A@
NP4+b7,T=FS6C_JLE:2NZG-GOe@<9GQJ(UL-<BS<8Z>c&2\D6#5@@_d8BaVU,DV]
S271:.4E3R3B=)8;RQ#2MfaI]QNQV\6-MLO5@4LF&\+1CX1P2aXGFK/^D)3&^F#Y
I/E0#/UB3b77:?/(4#0H)f3923KB+Z:N-/TF+S>g1#KUg1WL(C5HAK<bNf1Y<R^;
WEEVAecW^@DYd^XJ@JTBDG?(.[;g>JRM@RGY1.YX+Kb4<eD\&.9EbFKTLS+5^da]
b-&N(S4#?gefdZZfK/5=>ZBBJ/+-5+7:+M6KfeP>W5WIKN,IcB2QfbCg3P[c)<E.
Lf)Z1S4IKIN5)Te>?#=].b_VN2^/_6Za0>EdN+J-Q2+GFL9Y3)3+e;8&;-#cK.M=
ZVf,/RLVFFJPE06#&D4;5ZV+)/),O(^F+AX-0;9b.T>T[C_9g]bFW:cO/+Sd4>]5
[^D2SQ_E0;6\P;bfIS>JEBK:f[^076]4#[#e;MJT@fA.JO@bJ(K/NW.9E7ERDJbf
8:<5D2>G]R&)fBC25,42dM7-7V=3N+@d4&79XG9d[K9860<3A+J8JQ?5Z4L&:Pf[
HN-S2VbD_0;3WV,Q#RH;(JD-0MgCP&#<W@L0_f-eF4Od24fJ1bJ3T9I1NTHRX@5K
BTeV&#ZWAIF6TVU7NgF106C_]fQ>IK7/HRR?-)I[B.f8Qb[dHQ8H=Z(F.5ae[g?1
2-B-4(OPa#+MHN0?BSRCP8^7ae9CO@S,&7X;5_Q5?fV\LEP37M_2b6C[#YWA1c.d
Hb>.,]aZ0@)IQRNOK=Jb/R;1I;;NQ1Z:HG&c?J?:-a^<2Xe8\S]RfF9RYT[ZbY;=
(UPTT;]N[dJE:2Q#e_O],Y)^[+C0^T]2X^A(Q@TR27+FI)_W#UF^(S+)ceQW_8NE
PDW0^C.\XK:,Me+GM2/>),-Bd(?]EVUQYDO]M+.-:-S&C4(1BZ^[\DL=JBfaQO5d
4(]gMZSEOZ^B@6WHOfOUK6X(0BabbVc4aCLG)2bZU;adQ(a&,P@(WE[E@)ZI[=TI
WCYT)dG<L]J@_Ld[:<d\e+3D492_ZNX&^RFd[N0#b9eK<f?P8H\dJe.L[G^\,9fa
=]U<NXM.NPS;[-25//g2<1e;W&#FP8+:EIB@QO]c<-L#VDNe7fQ>eY1G@bb2B(NV
eRECKH^OSaOMbgbZfa8He2>OGaY;LW..dU57.CF(:>P)Q;1\B+E)\_7TR6230e3#
-XMXJS\8Q9R._X9WbQ)V\&\fgQTbb_<@45@94?Y6N.9#LZYK_U7P(U/HB,_54a3K
EeZDU^I6A+5L_R7.#+HMb=AXY<MJ>V&XM3CfB&0g</(X1:1bd?1:[N./\Z=2\U#.
dAe.:eK<\5BOUJDf-T]g^^L=b8^/5MJ+ASGgR)_C4M;.JB3/EOLK#b9BgePH4).0
Nd_T?6;VPL09GE@8>2e79O(]QHX>gW?W;^)7>V7B-a(A5)CI1EX:IZFTT\\^OPR=
.?-&5@W/L.H=T0^b2]-51Ed6;)&]-5B#/-Z\8H8g,_T_N,AO(71CCgCYMRMWW6E#
\\V,NS024&ICg^S[cNSc7>:=_0HCFDDIZ(B]+M[>fTX2_SHX:#dTUE)7eRHT]cPY
_6G=^53T4Lf5)A.d0):C2=\-HNTQQQ3I]WCdC>g00>\dLK>YAIc9?3GWT:I6BBXc
1gd=80faQ)W/g<5HAL=SAg83<2FF;>3A8Y)&6UEQ;#LA-N4eH08QgHWfcA(.a8[a
c?6D=H(N7Z(/Z2@(aLW?]IgfJ<A7M_CSQJOSUT\Z.X)YeGae4-gdeUY)/F;XTBXO
O<@2?Cf<=?\XJK?>(YMcga5LL=B4\Dca)Q^^gda@<eg,D52U:^bfCeb#PaeK&@B)
/KW^5_aT:eU4H+,f2SGQ=UBb0Y>a3Y2SU-Ab:7R8^QW]P<JC54Zdb87UATE=8_W6
P]2:#UEQF[.g,EVY@Y>Q.g4MK)+G]B5J,6W(XU@W=@e=CF,b]JPYU1Id,7\(&KS)
C(M]N=Z10dD_IJPgX&TL.RMK>gcWa^U</3QcJ#R9C]\19<,#eYSQ@eUSB#e=?F@:
YX4+4>&\ID0[\1YUSO-<3ZfO@)K#bG.?d;24E-II:Pe2PCCPLJ>b-:&P-EdZCATe
g))W7;[&-#A/?+N1?-]bBVY(K2UcC#@,O;GFTK63V&TA^TgU^-HAF\ES8]LNOZ+L
bS;Z8=<E:J+);ZI1.E)LffZ4<I)7W+fPFc[8.C<[\:_JAge2]U4-)=NG]D;W+-:#
>CQ3.I4d2;^SO=0WO/4@?eCf8fGIJZgY<^O3;e6T8J.;Q]XAVJ/1TK_GHYYZ?47N
J;fVI?2BV\c-ZH,Ga3_)F_:.1KU=S;Nf5<RC.O/HVKgO;AKFTD0WG^+LC@]MeGP=
?7>G:/g558LJQ2a<bBTCZdE[RDYRKI]1)RJ(I[1_;1)P=?cKWFb7M,HA^a#Z6=)C
(;6d[X[]S#Z3EA=NP-8?fV_=fM<YF3HA/a>FG[+5^[6bKGJMcH6&-5IM_Oe;b;?2
ER63?H;b3G?FN:]U(-PHS)bac^I7YcHDOOSVZ0?,?GBfcF7XgeAH7)6/U/L^Wgf(
]C.86JeZ?NF^;H^eJ..B]I#Qg?7-?3/bbOJOeDL8gAB9J?e7#S0.eY<H9)\9c>]=
9W@/RUC37Q?eYP_7];bTU<>T]VMD5<VPGf?M<[8\+HXF&A=QOAY1ae.V3))c]_Z8
bb3a8RN@&MXH:7+Q@W[\:CcdZN.OHB&4=.0^6PdNZ4^4#9)/#S5^8L738B+A9RI8
>T^[C<A)JfHIg:4P_1M?ScGc0b^a177XNgR1VOcJRc/M5->H=+&f1[<eYL_A1gB^
,V4>MP&4bS:MEfcgA?I)Ha#QL+:cVEa,SUYL&d/5Od8aAY=YF@^]#JXK1RJ-?M=S
6Z.=C9[1.H-BF23J.;eE1AB.a8VeD88B]KD6BDS>T&cIH[Lg(@D>f8-/?=Hg_L@SR$
`endprotected
