`ifdef RTL
    `define CYCLE_TIME 10.0
`endif
`ifdef GATE
    `define CYCLE_TIME 10.0
`endif

module PATTERN(
    // Output signals
    clk,
	rst_n,
	in_valid,
    in_data, 
	in_mode,
    // Input signals
    out_valid, 
	out_data
);


`protected
^5\c<ef#L\PF-:CX_J1XPc3O9],^9BgSFa)E)#I#4L2G(_4_WHQ4+)E1LDf:H5bD
#Q8ALX.Q5@Q.]HO8eUe(X27Ka(YDWaBU35=N:?X:3SRMCY_DFf9U1?TT,bNJIJLY
VJIe-F=AUOC@EB)b7_U_c[4A]G;#,:U\AOW,9Sf=P,MM<2NVHC9MDK_cFe(3RS,T
-3F<UM]<6FGW-KYGNQP(3X4A5$
`endprotected
output reg clk, rst_n, in_valid;
output reg [8:0] in_mode;
output reg [14:0] in_data;

input out_valid;
input [206:0] out_data;


`protected
O8gF-Z6NDMJF(X#f6PCUIU#QUE0\44\8B<96aME0&&>(+R3A^4VV2)c^^?J9S,71
/PD(;/8_C[^Ia?<2g@f.KAX9.U0#Z<PAH+X:XZH_Y00X,K&BF<]6d(MY5Vc=0UV-
2V@(_McNd-=SIH:@N768AZ-KU,YZAZT&-SXRL;daN\YF=b\K_O(L9?R_+04:HG4X
ZfD=cS;L]7RR2M.PJ#.b(2BCDSgdFQd5?&<EUdU#W&4:1>?AE16(48K.D4LOY4^^
#77)>=R0V9Y](2&N<0(XaZ3Qa=8?-6^W7cAeM>g8E47-1gg[\_:W\B\f?5DD:DCc
e7A(ZP(eQS2H[SGa5aMCcE_:+fKS.56e8W&.U7Z07fJW(IUYc5:G&;(OU?J>Qd2:
OF>Rc<3gNF]d2WV5E_gU<H+f3RaF-^Ee?OIXK)E?RH#9EGfAL?W420>K-6D+6I?U
1gefY=@>-5+/&d6#Pd3#/b5/#9F^MfKeT.S8BDT77M)W./INJR9]/Ba-7B[fbPX6
MK3T:LFR[UW(+@:=NK-<3E;]f6\@=-_QG&B+aHS2F:1^@IYX=FG==<d+e@/:dOBd
N/6V8UY5RN9@V;&21^.;A5K]PCbN,CL2S:/ZV0]X(Q>7J-:#;bH]BfT&4VVVG3&O
a6GVfPJV1eCU:</]\89Lf4DAR@J@N@MCe7K08SdRV^KUXa7?&;cTXe4^IWNF/(7f
34g4/#4LQ^Ye/^@fP+4NF^CFJ:8>2CBD01:=]GKbF.HPPg62>_@47^@f5d2;]R[X
9e[cMS(0B7Y-\#WdV#HC7+U#O]2H1-1IP9?g&-^&R6TO[O@cH27X(AORHbeD_FLW
.6#;C;d#GU4[&FebgVWM=;1F&23<XK2O0:1GfUJf4=:(P?BSc1+:SZ<ODMG2]D4<
,2;B0;<3&g;8;)(FL)d>-3[;&bf#4XYA=I_YT>ePP06QdGWN)4_cZHd[K+UT5VA(
FPFLW8[gU+gGb3H?=5&gR&^=AdYAU:<YDKJ1EQD:.XF&?c8TUe#Gf.MePC]KZY@e
RMM<+VI2);2R(&UR1C#BA_a(_LFc^TfSbdN-fS@,@8E]BdWV(a^,5&X3&@_&>+IW
eA\4);eU?C/a+BPGf]C4b##f/R:dTT4(RWe.?/O6OUE;f[>^TK(.,7M-41,MF1:g
U=YRSEU5FYO@4J:0X<fb(9_(>2L#^9Fe7L7]X=+6P?BDNCE#f>&0^HAEB8Q7WM\X
;Q4AbUK/+EMSB\(MbePgU)1S@[&fd0cdL^JOQUb(Zfb@E;IHdMHcN(F?NBTFS6.#
2?16#L+@R98FE-0[W;D1Z)I)I8bXg[#d1SH.2)\(^M25FLYO/M[&7PTCWCMbgLFY
4:_)Y<3E0KFNJaAg[H[.TE@9,J7CH;O=g\3>3R3]61O8eT(6Ae7@_RYH.R:IM+^]
QBZb?NI35A8Ia8HfW=?UNZ#5::XMM4HLHcd)bK>-BY-c&K>ZN_T@dP8cQc0K=;7=
6?O^;5E3LQ-AQ_@b2-SLW.70W>P7TJ.;>.5?\7G0[1:4JHY+D0F0?3e:JS,[Xg9C
Y^5A.SI8/24,^JL>dIdB\^I<556=#();P[Ye1TL\d#e12.PZ-b[]J0f6CG1DUPHf
94P.;(;SM@Af=eLfOT=OB27M16.d.<0,0:.8A[a]WA##I+SLF+77L7@?LbJ:g/fD
YT7S27?U(?=EPda^Ad/96<aRdNI#XRDD@J/Fd&a-:eQ7L1W48I[7@Q\G(OJg-YIM
K>AcQa;R4T?XdGdTO\C\9J.K&HVd646(JS&[YQbJ#&I5fIFG>LH99:RL=YVE.gVY
;M6E3MSKGd\<8;9Q.^TWG,RUI69E1V,CP5=D)>a]b/=,J_&S3dR2I6_L0Y5D7LH#
e38SgGBVRb1Zd>-PO;SGf#>/GcF3P8d:,7FVAdE<C5?253Vg_[e\B.HV>7F_1;Z0
B\[OY?fIeR1)Y(c^T5(2N2LQ@^TTSCFfJf)AI_4H&F+LDQe97&eEV<GA_QC#YG]B
AUd^.6S&W8)Pc1L>MW&eLMUdH/R7\,(;@JQL8b\+3HI3W&K.e^<&&I79L.E>O=C#
P-UYaWC906DA><L[4IaWdNALfe5NgGO/OIZ[/E^U=8G3_1VC;(-V])^HH&ZICTeQ
;5RE,f5&K>08,TFXOZfX\<YFZ_,9B?9-EaX:N6(aV&@3NV8TFKRJf0AT<7HLL;G:
?7D8][3Y/M?RT@YFYBN5B.HT:3+2T<g\-N(@-T1,;.ZWgI\0HD4Qc>gDf-O[UQC&
/3PW((MgE.d#A13#ecZa6B&9g\Ee^Z@6E01C4@T2.ZRG>/_(9.Lf9T>g;&N1Ud^7
d?2QE;@6B2D@I.GQW^@?<fH(7V\DG=J[J-17=A9:FA?/1C9/R;J?fd0g[aCR>.#H
EZTOf#8SHNb@?Z][^[M3^OKT9e_5a7g7QcG[-WB(Wc+7U<ZbgC&RVM-;(0[NVZQP
EZRMNK>fgH?;L7[.1@6S#AFVb6M2KA]:2fYWP/C&[bMD?T?@+800X8#d;-Pc^0^K
O)YUZ/MWK.WJFURWd6a&R,6XJI)GM,7_-E7DV@&))+8BN/XOW2U5B0JYg<^DUD;I
eLFbLBcL#fbc4_7IP,Y&S9cLaA+YYKg;UMcIa=_63LbW_^6cb;\ae&eM,&UA[c_Z
5&c9YF007/5LMMbF<G=R4=OYcE-0N]E4P1J/^/G5=Cf3EBPP9CGD0;gRZO@O.\0e
B2&DK\09cX+V/gP+>cdS42H6aKRJ7ZUHRXQ10(8=bRH([g?OaS#2U(a@<>M6BR[=
)[\XLU=/8T7TIF(a37(ZKf.)a:g9c:bD0^&(T4]59&C+:+S9R[G7]egg2Eb/YVK,
Ad_1-(I:OKc5_L[aFcH=Og0+I6P&6WX:=.)@,J_cgP4MF-KVQ4M68^GM&8(3L6C6
O;c]/>/ZMF4-)gX-#/L>S:)#5NOe+b^YJ@1_;I#6K.THaFLJLc)TL3N<[aVJ\6OG
O9<O_@2BH8aPP7,[REg+gCf2BK#1]8C#P0B1TO6(@E7)HdD\@7TVK?\YJUe,b10Q
L?ddG2QVXO&O?9V9IV@_+&BH1cDO]B[3ZR22)eDWZHCTQ7Q[V>8#-ZB>JP52Z#^]
.\K+BV?8HPO>0d8e/d4=W&IG5[e].1&#R8^b&T/b^XbbZ[ZcU@(OLg:d<?dO.-?)
,/H?a,JY:NR8#;-0cZNK-eI/QF6747,WD4P[00]I;F(A:+N[,HfEa(EKY\.)ag@&
)1C..A@_+P=262Z.G[f+aU@/&=DE?:Q6.^aIUeGg+TD,ML^-(^QK\:/1)JZD^O4O
Nb6X>S=LG79I>@A_0HTLB@a\BE#VM8_V+8KMM1\CW80GU@J=;Q2[[cID[bM&1^aJ
]73X)F]U]e<P##R?1/[5OD5P5QWHO9N1TgRJIA[<VPSQJX#._e=8]5>:>DKJ[HOO
)<GCD)f0:P4/M>0XAbB5BTa2f37/P@]F7f,@XF2^0OV/NZbJ=bbW(FN&GHBP8)VP
2;aR0<[R5cNX[CLY/&G\KX+OA7SO5e&;&:N\+-Ce&Y7dXAIe=J=RY-G@_;^,K[P:
PH7ZA:&a<<VS_Z7;[.)_OJ_VXMUD6LMX?IB<3&Id&eI8F1M.-+E+Kf.^Df_:5,\a
R3da)?^6.LL.XdWOHeYT&=;=N8X-NGXV?gOCN(BJg,GGa(W.H?[BCN^^=E6S,;8Z
bXcD>-H2\R>^9F2ZM&7bE64+6F1\/.-U#-1X]6feAPBRdQ[RNVW))cE,d(O]fW(B
_6RT3Q557/=TLYRJA9G8]2A+K+54L(VR351I5)SVG[=@DBMDZG+\]\0(,7[-(GNV
]ccH-==d@6BU91.OB(a2Z>N6)XO>)Kd()N@4D?Cc:X<D:PVJE(AGe6WK7B4,eY2b
cH-5Wb(AFO9SSM5d=RRSLOGb](ANOIFe#LDP/a.2=@=\;H75L]TKU(#+QI=2Qe]]
^SPe8dCIYE1].\UG_Y#NFL@ZV[d.7dQ>@V3=MBF.E2J9Bg5f0J+),fbWD08U.1^Y
CM=@I.6>cC8_]Vba9UPAG3_0,KB<1/[O29W=KacEI.?#g#0)XOM[=e9HcLP0K2aI
Od<AQX^Vad(9,\9E:KB8c4K:P=4^:^eR@ff]OD,BI>9VF9Vd<&)4?Q?>NW&dP[&]
OJY66;\\(8c=]X\;&0F]^_?Jf+P<JX;<+HM,VYc;Aa+ZM(eGU<CXb-a2J_.cMG8V
BKA]WH#]P<b))Q/<U\D.]11A.6QEPK:>DCZ@#LfXYX97&O13]YIbV4^8&P?5T^^>
(9?K&[I-9G1)&cQ.\/==XXRZ0W_=RB#9ERAKdH(bX]?f^O[<<GS>)IgY,CM[&.G>
EA6.:(g>ELH)Ob9XaOD-74Y,SdTMZUE[JJY)O_?:e:2\UK-W:3CZb=WU(ZXM4T59
\@QQ3d.M2cOa[CK)E[f9P-S\X]XB38=^N:K13_gI-V_R5PN7GBG\b.PM#),>Kc84
+4#KJeHMWNM>^K>/W,T_X[W?CJ3(Q-a\V.(XQM&1]GfDSBWc,YS4R>Y_T(Y@IG<>
TLM5M1QeV:.9(<^9M)e6UGQ+A8#e4RKbN5NTK9;?.@KV<C[[IR43+8U[Vc3R.:NT
UY&]WKCT6;9L7QDBF=Ne]:cP=b+3&H?#,cAHa>aDS7:(NLg4d14F34E([_Zf3J+L
C_:FgQE]J)KdIUb1^<S[-F<;@T[2]fXgd48gG<MXCAbH2)6Z>.8<1E\H.P1EXd-Y
)fG_dZKA/6Od3F39[>R\/0?[J_Z<,>GG?+a5-gfOb7e=+a^)H]=;(Z2D3gMOE+L,
5C=VfU#2+AJ:MC4cfRL^14P&#7Q[5X6.P7,_NV@H=QR6NWc@:/4B]Yg6c=C3]_gc
Ld/2+gVG=Z/PeT2,/M<Q_WGUCY)+@^QX@AN@#P1c@KY;B6-]QVU=dS.:?g.,f_7B
fZJN[6T\8VbS5aOgP&VW+04:KbSL1c7M-TTSRR)f<CRI_]g.-><@1#YU131b2DX&
UYTXH@3VAUaR3,fUCA>\O,)\fZ:R]8H4]1Z3EKg?NcR<Oa)V7+<]_ZG]b7[-Z545
b]DQQM;c-U8N\H.9E,;C^<3DCW;(XW9cfD^1RX>1(EJ+U(8V=ZWR-G/Ha,#PJaJL
IOAa2U(@e?DJcg-5UMNKU/UY]ZNA#_?ZP\W6;/XN9Ld_V4O[J(:1/TLe5.:>/DY9
G,e)U+YGW_P<B@CX8NO(10;cEC4\6RLaSVE8:aT,ZH5=UX.TZ^KYUcHUHcA2;LMV
>U;9c-[fB656a?W,SR):.>ME6HXB4V#(_3<2#3=@[\)QD04#WPHV(EH<W&0b7Id@
+P)>LG]fJ31^,bf>U]/c^HY27@eI^9Tdc+5_a+:?b.f)<H9V9a?&fR89P652G3HJ
XM#RVP:VZA@DYdRR_;6IN_RN\+f8->MZ#PXdSaCeP\[-]0T63c?)L_SS<\RMU,WU
&3HKeM)gKA+7VAgdB,3O7+AT\(@PA:B[FD#Vf0GL1SKg)CPfcC;\->DIL^_S;dQ3
L_b7NK<A;3S&KCa9K[#W4Rf-bL;QUCSMa@HXbN7#ZAS4JHfFHDgATBH]#&F8b;8;
S9U3-gNMbNI6^8SG@.E0OfOZ30RGb,X:_)\:,4I,FdYEbOGX(0T@<UE#FU8bT.BI
eK6<fc4aRC[J@Y,2X^G_:6-7HN#HB6A\^B9&,)GE-PbA,gZgbP\UKXM,KLSS@U]5
@O<6W1+O/8A^BfP3:FR7Y=2(#&Y918+?ZCA(E)Cgg^)+Uc-ET4&NRc53GZ7YYP8[
H1M+MQT&\N[ZMQ?M?1]U:/+G\(g.&LDX7:Zd4N(1b^ecRX)]=C;>)?=eaS(U&K8N
f72HdV>W#5[M\G8=VYR,CE87NE?>c//249)dPRbDW8SO7L=EPeRbP)/E.+A&KUJW
EBM;CF_Fg:UZ&AX_E]TfD_C58e;?63NR,:36Mc<5&_IVTYDa6;.VP0/))@>D@I[S
GQa2_/_/AfMOEOFB0I-RZ#S:BF5HU/O.9Ff,?gJK99;J2P()?8U)]fD#TQ5=NV#T
4L1)>TNND9=PIWL/E4aO6(1d43U3LfR5KP32O^(4;D>M]1PI.?#Z?Q>##]TIM(fN
>+#ZgLD#S[.E<N)Q6_^g0+V-A&Q6U#Z+NF/Rb3fW)&-,Xg7HOVE&D+(fW,N@B8c1
&P\g8=1B6e+>L64EP=(bPD#H(#bQ:I.[Re@(<S@Ue3KX-\;b</a.>9#^\X;?,(F3
8\e2__G5M/[8W,R+@gf^,=C+)1OD3WHHLZDH,(V;0V:37VB2AK><G03Y@2F&]]G]
2+T77^<e5CN64Y#e#/AR6A25E4Z9GZ05W[TW>7bG.Ma]((2R2;P2VSFcF#YE9a0(
+A0>Q?aZW]NN/)<#=e4;2Q>2PfW.GKA<W7J,C>b,V,KKHQB6fWbMYOdHb<2P[Oc;
\L0<NN6#^OJ3L<f-2G:6@LAOM/QgAX=62N(C)E56:Mc&M;.#,-V.b2(80.,6<N)7
G4g[9a#F1[fF=0)<,@Z&Z2YLe3)U8I6MATU3c6Ge_B3W?\+.eE5a_@3P;:I;X=9I
d[.=:>4BO@GV2([)5CdHC;#O<?IWZ2STRW;9b(/f=JDa:M\d6&IA]P<_J8g8?O(_
e&@469=S.+&^a#(-=@I5O.9.bDaXS_(e^9IW0F;>[&MX50c&IGeOX^e?Y:LXM,DZ
&;5Jg,_QbJFVUJBH9#HF@bS)MGHcWga-HPW_RGB)f2A6M#,WBHG)Q.Z5L/(OWB^=
^IUfRKO0<R46V:FB\:K@ONHXWZ#TG2J]:AS,R3Y4/UPdae7W@;26IgZHT<KgDZH&
@#G(H+^8:@VbJU?(#CZA/].(_QFKbb<1@V.W@R0Y_4KP5?(0S2\bPXCO7FB:AdP]
XXNOFHT70,AEK[NBWE-N+-BPI0E-G&L[HNb0IGG(#W?MD)@[8\75F113Rg=9P0?b
d90W223+CFPSRW)>gW=\[W=/PKgb]/bcF-28A8Y7X[BD)+^SKdS8e<e.+2B\+J,[
TA7##e+[UVd+3T8_\DQ93)#Ng@=IGe\Z]WHHTI;E<4&Y<0PC>P&./+WVd2+,Va[J
AO_])BKBf]f;EQb#S=K<Y2F9_UdaeAePaR+5KP03U>Jgec\/XK1cbEP&MOa[-D<B
T=g4Z9?FVPL])SSbe3H3GaK\7@C8G4^V:,dL]IDJc/3.fKg@P@BDRNMWdd#e=R#,
#,1fXVAT\&:99[(cO^+CY4:\Z<:M4?21IJ<c[7MV4Z?7BKFK)..C^SORUNU[DZ0H
?gG3TPAT=2dBK/>RZE_5:#U-\F_Xc:B6d,YagG323?K1#)XAGA#?6Hd&FG.\];YY
EQ\GD+WD=YL47CZ5UR/@3@SY-+&(8\^N4_N,8fV>:S]&gJKOWXML0+JK)3^85IM^
JPKa,g,/G[TF_EG-8O-GDZd,1:EQe8G2EN;=D7Z[STZ5X,YWf46X8DGHY^_[1DYZ
C@,gG1e80df9HQTa/(GVK][:T+\U88bFdcc<_PU.&gLFLJYbb<P]NF^IT#.ENReS
.>38Kdg?4_Ke^1&=[8)HV,]7b0>C,WQaTY0WHPGIN3fe4C56L:dJ-5?/Ua8,-K]=
aWYRcPP=^3C2=0g7H:b3JTY@L]Q;FTE/,eXC+>R:H^??<]N<f5+b-3cF.OP]GfeR
MTB1GVXE98;#FDDX@+])5EWS6(-[E8E5Od@?X6STXNU/^:;VO3PZM8V1=[g3U+8G
A&T>^3JfGNWX1XbH,CFL:Pc90dg5;-BDBU0LC2__(=?O:a;(XRO:\0UgW&SW7FSY
(\7S=7B@M_AGf=9L4(H_Vf[]OI,DNUHe0KYe/3YK5@A6ZXc_eGT7)QR6Y]NG4C3G
(G:2?RYFR=YTg?;)L6_-NE+O[/#beBG>?EW^fG8C8SQ=UWQX\+F..a7&1AaJYcNH
5bX/K)199B[A3L+L^HaSQ5Fe_2MKEe:[eg_EbF)Q_YP]D+HSD,[UH?QZME=NSYZ+
ecPEOIDB=[1S-QQG\FV#:RIKCA.S_[Y>Xcf<IHU/b4<ag0]AM\V5R<H57;>]>d)U
-E(Ve5(aQB.9FNMJL[R1F+\+GaO@I.NVdf;9,&];8QX/.BL13(10L_.Z6S@>#gBO
[X;DZL5_d;2P&DcB^,U#>(R4W,(P[_?V[=CD6(DZ,e3CH)/@UF>cg=+7EfK-Bcd@
@XR,g?/0,BQJ<J-gfX_A;<[YL=\@,C2+++XNWVN:@T66?F]g?>02g@RD>9IfFS4E
SP)8NZf<MNV?D#L4=W-8\=>H2Z]6,W0UWHFA^2+gV#N>+1UVD2UU+e0_>>LOd@C#
4/B1B:WBS5Ddd5-A;0,;&cE]CM]==;N3ZV-EQAaIU>6H?B4.G^[@b(<4UT9cB0&D
ET14bN?O?4P2_f(UJf3AOE=@-g8fdI;Wa]__=RVfT9,@33_PW7DN3aVQ3]6\^\/Y
M=U+MHN2(BTLLW2G^gA8CK#1=]Y&9.Xe^eTOeL&XDYX@(CW,:<\\9^Z8F@&#FA1P
0S?@A(3,)R<LHMdS8/b4E)#EdO#Q5P1dIQXX;S<(HX4\66a(XP2QeIG+^M8c3[[,
b^#\)baA=Q.#@+VPQ&&fJ;WVN#E(VKa7BcQ8ReX+H&6LP3WPF[MDHG;;M\SDI#PV
\X@U;Xb\HB7f9F),OEU)g@d&D=0T#e[2@PN<J5T+8HPQ4>[<g6^&TU#bI6>Baf0H
Sd6)<EKV1?:KOe1EO@PHc70PEPIA17gV_1ge82A3Ub09bB>^CSGN?b)DJAKc_.e-
fdf0S3:5W)#_f(gVbDM<bM/fZ#6\&;1KD<)(C;22ZcC2829^\-5LFH0#HK<M]faF
31?,=d[ITF0@R\d8MVH]\H@(&GK6VJ,TD0dgW<(cFKZR<+YPA94T9HKCd?=^RX/S
#TJgNNBg5AMLT#P^QK<3#7gQ@H5CM/=WHH)5T;5e];c(Q>/:FE5Rc6SEN0T;Z+R5
S8(;Z,,4[79/Q2-#D.=REgY+MI@QDDDVM6:aU9X9SN\RGdZ6N3f20V-+VcYJ<8#L
MFX9aF;]81b\HKN_2^:d6]g7&4&8TPT<O_Y:5O/>R:PQTBfSac6]7GB16\^T@:e#
[)-A8:a7928H+@Sa>Y.gQ5;OYZ&df#P<_8dE>LcQafF=FG5B<PgL-bQ3\@\e(U)&
;2E.CJad8g:O=f(XJ4aT3J&gc,=4Xg:KH6LBL+H>_e9:fCVMaY_A-NLW^1&WeO\W
g+JJ&H2]>7Lc4PKS;FXRF,&R+\6)Bd:]3XAK8<XSPIYWEB>D(XD75E=.2WgXR2X1
[H)-+d<XY28B7_S_02;K]&;OH9bWJ#=8AcZCaaVSXBEgXbPDP3ZP8R@>X^VUY>:X
g4N84X+7G86J4=Dc8dedMG^.;cK6Gc)UW;K\-2R=8;>4gX]?_:ZA/HZ,66M<B(1<
5>fL]3S8GUA##F,]3>K:EQ12J_)TDNe5f,XGd_GaW>Df&5#4RRb,8>](VJJ,9DQ8
Q;A2aK]2A&J+]0.b.[.5aWH50;A23E2=56_?NS6G_/<R0#)X#1-V-a/#YI1E,7JQ
SHGQ)GA:CBKfTPC>Y^gPX>6VV=.XN/Rd,:g\Ff+Z64ERZ:dH(9f>?Df3Y.dW.dUa
E.cWbKXMceLF(+386Z8^]>>WZ.8fTSfXN66NN:WG\>\X<+:IZA_-L@3.QBa\JWCZ
&;Db@W]TYcL8&e9AHZF2B99f^2+f@XfgIJg=e0(0Z5J2@:QMKQRWf&SVa.?VgHTA
;FT,ba6=O1:BgU1F^7e3-[L[AfDQcZf#Z.]6R,-8S&YaFA8/MXYMdZ-,E8EW)a-F
aZC,fD/,;Yf;(dLHAQ,:T3:H,W+Q&Pdc3T>2)c04SRHU]fJeY@R4NeQ,#-M_,G0g
_;&8-3e&YG=Rb)c@EK5^OT]SB+-@4)Uf:G)9L5>R2(+LZ5:ST?S0<aE\2P4(ZcMX
C:1Ka2==_b]ZRe9_f9:U#Zeb.1c_Mc^#-aR[20=UY(cT&bY01^B(2d7[)1/QZAO2
Tgf7[J0\&6OaPBW<a2.5=0]CY3g\6<L3#Zg^NF/G]AO5QX]7FP^J+Y1d_6g5QGYE
TGDRGCL5YE>.8L(Sa5@6,a:\V/^/=L87NcIW5K,^</D])7cVb3fDbZaTE4VR?bX/
cJ=^G[f))Y5>I;8@]<e(&VEOac/O_1EH:Q.VVfaNEaWdg#1NOP69+Yb[35V8g[8X
.0,f9gWFQ#(<X-J+A:U^BEF(Wd@.Ue4:,?#Hb)=F4fbU]3S=MF81SIb:Y>=G-cfX
FRDNg&D)99e?O0[A_T#4QIgZ=GbSD)GR<&&.8]T)e:((M8C>a+0YceO/4]VC>.2:
@<V.e6>S,<=a^;c8\V,eINLVJA)H8.\6Q#X/EL(^AOS(X3)-YfE?].]NYA&caLM5
N.KP4c?c&-UC/S)MdUR:W09VA7;V.ZHW7bT#eU2FZ[Z/+,-UJZCDVgFeDKKO/K<A
7O;W?e//-FfBa-B?EBE14eN#f_2AD878+W?^5#OZd@QP-UL]9QL\^F68>(VM0((/
Z::fR78R7L2EFL[VZWSWLADI.-d@bDW]YD;_\X+dP,\Q:<7_YdSeS,Mb7Cd\-&JU
TAM3]#/4(8aNgd#7A0XEL\2TNLU]YbgH;:KGDRVLDUbK_K)1DF/dH>89]=#]0RgZ
1DV=F52#.bEVAVM&NL8H<QTA7\6a8[N3HC5\TAIT2\_S3P0MWF\Q/+S7,/Tfb^6Z
;C.[g;^XIQZBe87+cB.E]aMC;X#dTZ0D>VOIc=^J4F(45?4HS#?.1Jb8^d)Q5Pa5
b-:Oc@5QdD\bSMOMNgIOZLfJ[O?IV>/fB^@c+Y&7-H3YN77<LGF9e](1c6YN2KL7
66U?e#.NJ&9a&OD165O(>WFg=5b;b,EGOWN#O:\7,?19ZW<QYNC=DIQ&Y(RIT;MA
C>V?8eg?]WYL64LecZF7N9?J:UC5b)]QE<[U?M7FUV]MW>4^@,0SF^1JA-->H-I>
D#2GDLE,3WfGE2)f4WDVW\T--g1UV,6aLK9F6g0b?S#Xa6ME.U2K8#O5;(e@9R0,
7f\FV;gOfS[fD0\-DgD[3^PQO=D7N^7c(^L0DL)CQYfYUa[T;Kg_gWcURT^@M>g@
\Ve@7Oe^QG@.HNY#>&@@ALGG5R\0Vf@e1?:<0UF[c3T&1agG@IK3[1U6+b>AWX>A
@)d_LPVc>3a_D3;X(Mg?Y)M+O;8]^1>cX7H1&9eL+YT2I86?E]S7eK0UBF7SHeS[
DTTM?,_<+O6SfT:,C9SFE.X^J;O>[61)BY3_g_c,-P/X=?&G0=O-e16(Hc7<J^^]
=QYLM62W\<ZHS(c\[KdJV,;A>c0.#XPGGfYV8MYJ.LY=5BF]0Ka9A]=g/[/38Q\F
ORZI4ZG]1E0RZ=;UO2Z0=7Q#[T3:FC?Z1I9+[?]J\<ERZJfR]0/<]2&X3)KSd^OB
/Y)^DU[HC@)a9+0+DT;@,6<D)MC-MJb]/Z<0]S6d<UK:9A?(>>aM=Y11b?FW_C#b
cX.3Z4d@Eda,)YD/.QWA@SI7S]3F1:6O92(VaB0NV=#3XBg8>37f=dgE=DIaBK:E
U8c/0.##9@A0aVTNI_9HPE(,-^ELYGW&#NXc9TFb<.;6WYH40;ZCV:3R7cVU(,F&
DFC#I6d_V5_HH74_LG^5A3c8F)58-Y5OK-[S.0JQV3T]c>E]NTfQfUU-ZFSUPYe8
b#QY)MTeN)V;N_#e9D<;Wa8&e:YHZYJ;Y^5;(X^6g0R7c8&:ZOg\7(gAd[SG\(+H
)0ac1gB3RY>HTb-ZPb9e=--dX8[911H?/<2b6P7Z=8D__e:@LegRM&-:J2[I+Nbe
g-5c-+c_cYBG0B7NVSUC87/J&AFQ/44ec/+WgY2S=&1^73IX:_4L22ZJCYR+VN2G
a5(.3IJP2Y,P/eW8=0\(E^be7X)?;8ZM#K41[UZ/L^8?6&WS8f,11<Q<f]_TVX.=
d2-J>fSZ[7-HOeB-ZSS=B#B&^Yc@71-[IXEU/_EZZ:\bXJ;4G]:b\]5KI]<U2R#(
W<H?I#9H;#?\G0F;6C_V7Y5<9HHYSNP+.FU9/@S8(f-.ASWI7_Y:&ccXIM=BMN9Y
5[5&@eCdbfIg,HRUI)4gLPWb\-dA6)5)TME\_7X#6R<c1eO5B:PUQ-E(C8-FHg[5
[Cde,fAU5](^E7FUSYeQg=<:FJL@[=:C@V-IMIE)&d#9-(EV.D@Z]Z.5];GKJBW@
(K@=+ZJeKWQ#APgJBf.;aTZ\^FKJBf>\ZWDR&0,T-,L>@gR=TK?CSZbNI3>5.7GY
^)K:FdEVG\E-NQdTV4:_1P@1gE:D426=(=Cef)-d4cE-T9XJ\K007VUaT2^-T3]6
>QcNM(AO([DKf#>OMd7g3(+I0M2d?=J38cAd7\Z@&#:f+V>L1KJOR5SeVJ1W;0O)
E/W24<I6#a@WM89WH#I[6C[-g/b71VT5NP#JC2Rg?cZMBOL3\=S>D.7^JFOA&:Q\
;[<KZCBQ.W,,EeaV\H#J5,=-=92Q66AOY6UO;\D?F^2QfdL/ZS:ANN<D&.d=,MR[
dM_)ZVKV1/F4&.1>H7)]EZUfU2NBeQPa8/\UU-TD+P?QMO&W:,--GU3&@X@gL6:3
Ce@g@&-Z__BO9e[815XWbLEd3ARDOW#1IJ_4.6_(<P)@A\GG&6VSR:AX3H?eX02;
/A>CWP7PJJ,gVO[V8CQ/g)egC,C(J[dB9W=(TIF+37/JU\D/;SI(_HWCS]Vd83TD
\/@aHKYL]TWP.&Z34K43Eb\9--\K<VIVa2I@Ke5)T>&L-FU,[B#1b?EZ-U<M@#Y2
3--TWL7+=#JCOQ1.^^+H>E.f3;][G()ebS1&19dY=N5GL1\(_<8XM8K95<]_d;K+
73,01ZObgGQ;/P#)5EFecf\V#T>;H8feKSQ-IbI>--EG-=RYK?Z31b=;;I7cb;R:
K-UG?5[0C?>6dA^HP/1,;Va@O]#A&5L<c7U7/?#4)7Sf&=EQR\[=4]TH0ABNMYEb
GP.+#&;)]I-(LR^9BUE.QI=3\Y]F8:QeH/H[+fg)]S>(gO90XK^)&YJaLg3,MfL^
+W;3Z;Dd9YRK>bccCRXf^UZ6Q(1R\Y&&B:P-.<gF=@5\e75c.WIUA2I6Y#_T5fE.
1X_Y0?UJ8DBT/#^-P5W;&9TM^N?H;6>KT71&NJ0-8B,6\,gG5fPbS[B&+fZY/W)b
-C:HSV0Jg/&07@-FORc=]^H^G?C,7TWY)c?bE596ADE]QW3R)[Z+GeWC4.EE\Vb<
R\4eDP/.1d0C_3Je@0,YG4,2Z4K[fO\OVX=YMNf#SXg4N1-81BWNZ\NJM>b(#Q:)
S+./W4K^J(8g#)X2(LPKR-fH,LaKLNM+X:F5F@8(g<9e+1P^D:,JNR,(XgIO9(Af
C-XT74a=ad0?&d\&]I^8QS4G@);W))<UV)_4XO\dLaa-Q_I:QW5J6?BJYNKUH&J;
UL;(,68@M=]2]D>Idfec-KY8X):CRCUL.>ZK\^1EWNbFF;O_RNHFf68S8VZNE(ZU
#-07UH;@4<L(S?^/.S_2]^-IeSD6)1R]c-S&,CLe\?3U@F8PP>f<GfII>a;aZ5Qc
;TFd\?cC&YPd(XDbL]UO?DET?DaI@:&(BQb^fWZG^.QReVBLH.&+:CWfg04/?UV@
;GY[cLW=agI+52=RG(FZ.eEVA0+?@+AdC1[Q8U53=GS+Y<IE#bLL0UB9fNU]#S?5
B1]94+[5d@&;HHFJ6O\,LgE#58\#[)I30ER(1TUa>=W]G[@I.WX>U[][ZeS=N0aP
Y>?_dG<7>_Rb)/9@FOX6-FO:3::-[EKCLJ_f,00QZ.PK[)04_CYT-B?0K2fdW<Rf
LZ[;&;>bZ0J.2_YK7:8c0ER@09d\]<#DRM+0??M2YN-E<YLVBWRV5(MgINEUVQ.,
/UgXa))4BCO&==V_\B<9(:EV\PDH[_S,5^<FNCDdC6.-:S>eRX/fY\QZ>;ARDVR6
,#/#Z<AMV3V?H<AY;<839AQO;2Nd55gB/MJY=F<9(&?49IIH#@\_-b:>HDB63>W2
1fTYH<a5\3ZDBFB/Z2YOH_9JUSHTAK[:O6Z?AU-VAP#A>V=)H&;c_BYS;Z6&Zc_P
<TUWcAf^c;DCR,KPNMK&&X1YMBXG>JRg;2cQ06fI4/g8ca4@8\[TJ9?^fAJD>>FY
YNT0::4N]?<Y[[O?_I4WFE<0JC@LPAb3[g.b3F;b/D8G0-WFW;((NAUe0\(TCP46
E;[b1[#/(TY.[X6PR=Tc5P3YQ>=8AU9+YIRHD?&UQ(T-6N[:V=8/+6J3:7(6bV][
g>CgF<+EJCYZ#_E^W;b(gQCgOK9G5M(B<GM(V]_Z17NcFKd=:GGE^EWTUK9=f).#
g?JVA41K4ZD,MNV)C^L>)SP8R/6#Y/0YdQ.Y6>Hc<-0C\?C?RHaWQJcSAEfC&5Mb
U[]^F2_@3>1gZ6EdP7J]<E<HH@X-&d=CU/DDI7IUdZ[I9\O9GX[RE:O>44=-AX:d
72UA9F/e^Z&L/X\@Cb/_S0+BUA7UR[.(H2HS2f(c_ddM1fbUaB<OVac1C@@dZ7;e
?:?.LK6/7bg2@eSa2]TAH4#&MXbgPFBV([L4(=#<92&-e79H6QK6ceHP:53a,,f&
)AGfS?A.?>G(\GI-@L_K]5K_&e_fP+TPFL33Kf3g#fFfed[)B;D+@D-TPB41e_Dc
I=Y<5;2J:^S)V5g/&:cP;d\>fVJSEB9_5HQ.E]?4UY,0FXUKB&c5X5Ed^fQX1D3O
K0\Jf,\MX3/MN=I>G2/YQUg=f(87>?RKL6TdL7+17?a9WESLG@3UBBB,>d9:Taa\
A&.5]:#>C0+5@.Je&5@GLf5PSL6^QTTL/=15Y7d2.RVXc5L=NLf@[&Lb1>9@\_:0
N4<U(.(X4.^[VQaNS9_7\c9BdSgY#Yc5&P@/3(R]JaMgHgH^5,<^GC8,OJS87I25
=/B>;;8T&0P?EO5U9LV9Sf8SGMbKSMCXFU^;4O;,c\,2.^)V??\/I#L+]>/QL/ZR
YIBFbd\^01EOeNgPaA4#e9B[80c02VPgR5.Bf1Mc07O66HbR:JT8ZC-IX=3+c-C(
\a)SIRAILMdHg_0D:^=WLVAH\?^KG[QXP<5E.d_(T98BQeP#Q8Y7--OGF3ERN\41
-:0/:B4>EB]AH&P<>=(P7]B2=),PbBOe=Y8&EgBM>9/FSMO@g0WC??[>1dDbNQAN
.egS-?>5.R4K:38aYA6Xd])_+cQU5g4B>&fG/;eP[)#DC6O3XHN,(,]TO.)+9U^]
KTQNW-E/d0=.Hg5O56Yf>c]P[/Kd9WTRV0C_\-OdL;-YeXLg7cfVQJZI2G_/(RC&
S<4)F6:26_V+c7Se\&I.CPOSWeH;C<895Gaa##DB&KAJTJBAb\-WeIVQL6:3Tac:
^3(X6AUIb2;;[&A:C0Gb>EBZSAgOVF1d.c&/C@+6)&1Qd/:NXU-^\YMOE6[\KNHE
0X,9@bFO(#d3=RTAMGe12L)ARF>GC32HNH@1^Z-BPOSf<2,7_>bE>QW)@YdG_&1;
;&=CYE2>Q25XHLTP>=[CAM77:gN1/1J1PePM5<&Zbe-9VCP;T;JQed8QSP-+5X?6
N^fE4&V8K@WP3.<JB[1adcGe_[KP\0c2D<+U/M6H\]NC+#F6SH?6d2JFN(PfM+#=
fC>>R,R_ZKP,,2_#6#E]/?fL8/PQ&]b,S8fJKG/#RSOP1A3b.T=f2Kd6c:,1LbUK
dbf@V#X3H:aY\).IB/<dcA,-WVITPe_f-::R-__[B(J,M57YVVa?/^9K30\.D(0O
@^&@fU@LZQYYG@6A[G5+I^R<_AN0<,9@G,Db?U0FVTYNc\1DOKN5B6a]]0BFL.S?
#A+TX?;.HVG4;GZ1PRK.>+bV:edcC2V@^Q+,[Nb[4:9Y0fdRC[<8bMS+SQI\?e[O
7I8]EKHBKYV2Z@61[BW[(LEcb^a7fA0WZ>.^CU0U;0.4UdF3RHZfNH#@Z?KG7c<K
@YIIP72I76#(-eNeYO0IPH49#aT)\#<0A4O_EUgXEAY)f6]+V3=O]d^QAGV7,9L#
6+OId\IaR9<:CAa_=,8I?f,D\,I^P-8G2GD=)><];(]5F?V4gXKWfSJ,cLObBN+N
e61A8TOK1FOGM(6F2Ge(/RIAe?XHUAD#6IB3P7gb6=g]Fg9MHcUL,Hb75T;\/5c+
4&U7MP@XRb@S^C3J-G)/O<^d/[g<aMSbQcM)X:N2a=F(6LNNETSf1VO3DJ3(4TeA
f(/d6MBMdT.,>D6]K_ILHgO_LeQ).de7J2&(#a^R-VVN]U)EO<0dHRXK#MWgK^KJ
\EZ/BYcEV:gI+H1I(93[8a;fF1<dOef^XZ/c&\]VW:W.6.,=gW\90HDeCbE_/1.;
1B2aA/gUVOJB>32)PP?/DZZ(5MP1&KRR@QPdV>G.DL:gTCKRf9PR#7=:UK4+OA9]
_=M,ZKX#(Pf3A@IGfWQ+6GRM<2)b3,.c?0a/.CZ4I>)=-83MGcG:RTS3_R((3AFa
f,[)d2WYVSU+1_AQJdISZOI6M5/IcVPb4gNcJeT&EYPOYJKcf<X@[XFe]VfUgb,C
0EdgN0^H\)1K25<;_+:JWHXD^Q[E67Kcf9I[KAW?/bJ5IA8/?@^4QYI@^V969E?5
C+,E+7P9&:)^,3)2bR98+Z:&SZ#IPa3-bS01.[X5Y68bg@2Q,@U.QEV2_K#B.11+
7&/a>]U>@]L+fSTCI-A.PV>]+[,?[93?,&LbLM-FND4GNG9Bcf2WLcDAX9\7d,9-
PG-GaG-HNZ)<\>FZ=5(>B?08/+.gHPS64S(;JQ>Q_RQ1?.(F?C\/FJA)WbW0Z,HG
5eD+-DZ_?#VdJgK?c.?I[1WgBMLg[F[JNRZWE5GDS\NW@51<CbN?bT?XKBM26CEO
(#RdSef0R[K0(WcVKL^SPD>6:Q/3K_1XNZ?Oc,#5A,I;ZLO]?H..(c)Q65U;YLE1
B+5eHgcY]9[J8Qd5=_g+,=;K3I-DH.][=gJ;9a#U:N)IGS.1[<)V-.=B3NL&Sa)V
]9-#+/+Mg\g(^I#>_KVZ(4K9W_^7_]DZW>W+acKJ&3:7&RQ#b(J3K=bb=CI2#G97
(0B4Y4=#0IDLLe++@;@7496_74\Bf614,KM59TGY/f7Z:B7g).1cW8T=GIH.]E>+
SVZ#2M=cLb(PWBUS@<D5YFZOIa].#aEUNU1R[,dFFf^>&S(H:+YR6/dAFTD89>7T
3\ADdfd3VL71[AcVLg&V#YF;3@7V6C:ceBEcg[8PIF6ER3)2MVO0eWDAYY_5#H2K
G[P1g#?YGLXdG_(eUcb9</XP_Lca^6OB:2EHL3<JOHCVP6MFbDX_=0CWNPC^:2/Y
D@@1^d]>R-Mb8PL;2c_ddV#/#Q:7DD1Y9bFgOSF;1?UfO__D14C-@=ZR75Mg@RW^
851L->c-/C)e&+ILP.JfW]4/E2O_D7(]dPZOWV7.<<:HCcfJ[]P(7g,NfcI^aRWR
LK.V?<V.Z,Ug:Ye5^Z_TUI_KK@O&&32_S.RH@7<R+/6N0WfHD/dLTgaJ/>#B1MZP
aL5:fULA\gKJf@;&<X+_:f7Ee=1Td,e<:KgI)?;-;>ESNL8W6+R9@@:#L=bXH;fG
-acagJcO>HHDIQ+[E2V<e/L_693DYIc-a#>/:QI0VIOV(3-FKYVHA(&)FIO.X8(&
_[d.(T>V,AcI_54H3BJTOP,&LIP7+8,GAY7@VE=a&-g76+CQbNZ5K4D#9A[NRe)&
.&ZJOBNf@d1I:f#W95IY.J9<a1HKZO/#5>2E3Uc[0V:J9Q-Z1daYS)<E.\RBN)1D
NMWZ<V>NP>.-:463Kd-7TAC4Ha=M09Mb##CE?/b<CE[T,Z3(H<g,0NTM.9H7E-NI
.b3<P4./K?HJX108<#R5USN>g?eT[=^XP0/^Bc>cAT(J_8)NOY3gZSCZ3]69OfeT
eD;TYAXE\f0YcUG&69I6(^-=#9)0)>Y,_RS;>O[GXa/WUBSYWc=6=A0B5#WH6,bM
0=YZWH8+[E;2J&=R2BP61a.Y[;,SUL5>YVJ6P_:>HFgTH+6aa?7#N-.A/ge(1_=8
)AdBdZP=eYf\UZ?+(d)-AJYFfbB-^dIFE;I8W9.GdWX5;VgZ^PdVUKOaUe81K0_Y
NY>+VP+4dN\<2gY]W7Z5ZbH5+Cc=D=7Q+;J3cgcg56/U]TZLfSgG.JeM/Y_-&U_S
0WGe6g<@/7/PGgg;#BJOf_563HgUDe<OH+KG],CL:<Za9e,)@>9SJ_FAUgA\X+V<
.d;HSJc\?@\3K,H=C?Rf\5BfV#>J5D\e4Wb7.)CW#_S1_agSRN?#5Hb,Q+e?KDa=
6c]U5H=dBC;K-#GRd0>YHCYSHJgI1@N(ZadQ@P5Q#46/X7SS^eNd?#T#@6b@;TJ5
OGNaI9aZ-Zb=NaYQZ4bIY>X#F1=4U)Q--\^FX)K[J]Cg37D)P-,e1?A^7SK=e]W.
ge[\Pf&WA@-A#C#7\=SdWBEda2eR<B;>>Bb)SJ3=,B]0J\Y+B3MXGU/,aOJB38SV
bHff1S<GF54GLS(FOWcF9,1AQ2Mg+WHD=@+LR2dHNJHPW_/T3SW>D>dMT0NZMg<)
cMD]F42U3Kd(BBP1,H>4T1@@A+R]^Q<O[[UWBD^J5G5@;D5J(Te;W.34B)Q9Vd[W
T13T2GN)1WA;K^Q(X3G,N?gf(V6:TM+d0LUaEEddR-,IS=ebYLd2GOOeC.:6gY5U
f/3\,I<=HQ/^252]\;fN5>aPH:gM;,?AE6;9K0B;Xd5.R-O]eQ6-YCY=S[GB_X6U
;.LZ#XS^EY?&QW9Q.]F@QHEW@:(;((aLe4<:&@OU0\RO,ef]N.,C3IWb<Y+U0F6?
D/Y\Z@BJ5)=1gb7\K?#3<8.g-d&B[YeT8X_@XGYK8?BY(_&7\]CGb6VU[^B)W@a[
O3THe?I:NY0KUJXH3F]@PZb6g^C>#b2K=TNO#R]S7P.Q12<I;Q<3LR-339P&;0=>
@G61+\J,7OWRVQ:X\5U;Y)B3).&?WT&K9S4E]&eZb<a]-AaCA1),K\E-Kf1<\F6>
Z7_-HK9XY-\BEU()4226&L7_K/[Ub3c9+fXbBE-&^#CgeUfMYD7f_cZABPQgLN[L
^Fg8]dATEe0g-LI(RCVd/CgAE>.C9.I:I]I+MPdTG7D)3NC9Z=:NA#K>BN233].Z
,L/R?f[\bFM#-JT&X9K1O8LC).SEYC2VNM4Q&(7/8K>]=L@N#6J-LOC5,D.3^;K_
WTKK7)5G1e-/H622HII=#+2-Ge>OgN,DL[8FF,0H7YFEL5Y.M+Z+5b:?.I6UE6SZ
F)10[BFJ9>D.EEY-ZOY2@f?/9KGS2Q_DYf(MOXSYHE1,P^PY<-#\U6:#/](5TF#b
E/-TaF(@5A<<I#gX7&(VJ6V(C;bTY\B^2[A+D91[-SI.+aOIF^495#g?M#K<6+O]
2)YK7_4(\?bc_W.2cL,^Y+[XCeM51<Z7U(7P_HgU_@Y4?Z9A-SfI8D\5ICd&TOGK
f9f/GME]ac58?B6&&ZMML)faWdR?4A>WG.?/HCTZ\PQ];@2<(30@V96?HA<_-,F9
WE5;WbPHW3Q;IbbdaQ#>V-=NG\F8@[^Q3=I3(\#,CG-NS>10MV.D[73W69(IMDH\
&&QIG9O=J23SW9/^\g8.9fffaOD^[59].9H(eTIBLAIFIK:9>Z.e;..H-3Ad6BU#
b#W7&YX;_L\J/e=Vf-Id?AdY#;@KM4CX6(]Jb<GF&N)3:D.aISPR\0.8SdT^@GMf
da+Jb^)K[X24RP,VS1=4CfQ+.MLWOJYQ<)&_3[?@B.eb=M0DgAGTe_f?\-=LBf)+
dG#:&.^=UZ@)Y_:HV,41E477T]T,G]F&&,_0?DDUS74BM36:_V--Jb&M@6>D;T2X
]]&H1:WR]0/&<IT0aRCO&XYg)_N-4;\fMLOHA7=XWg_O]XM9YP,>@,(X2gZ.5(6e
?0FPKF9cQ3BOT=(GYVC86T.AC.A_FG^Q6O4:>/4O#JGQTf+[b:R5KKgBB(IU^^&E
.,^GZ8@Z[I+<DMLB#Z6U,?TS+ED9;)4fXY/(39=];YM,F.W86.TT?QR:b21@Me/g
.B\1c>MA(<O/W+D_a-EP_W26.1;K\-/<:F:YFCMZFBLfK&FODV:=\DYJ=B.:cN1S
CZQY4:Z4HZQ1P?IXJW?(6VE;ZZEg?2;X)GJ;/I3c)V_>],?ZOU4=bZ]:?E#g0>SC
B:;cS=3FU&TG6M/+67Z#d7?UB^\f,Tc=^T_8)RNSCd_Q6fgU1I<QOLSLL7EGUU.[
R&6^XKR.3;)4Bf^OVAPI>@dcEgY.+5e0<I?P]e14b>2HEHa00Pcf252)eb:[Z]F@
-e(LT=CW]^Y]0)a[PZ#AHA(6VHQ3.Nc=3-^Ka^_EHf3<NXYDRe[MC6B7@96A-9#]
YATNKadcRaM77^1BVC9DRaI>Y&Z)&bU_-+;b3\35.Y&@QS:X@4F\#bF@&Dbf<-](
G4_^cO19O5GS+2aQ:@97gOeV6AZA+-F>JcDH?/K(cFK+fKID?FL-B]g&=a/-P:JR
I+94->b0HXHKI?.#KJ>D;;Ha40FBCWf5&&gb9.bDPP6>[QPM,08A\gW14#>0VaO\
CABM,V=1=C37bF8;T))IS_Ae]/SQ.U6]6eT\5c+c0I.XSI>?&-b[f1XI:g&;P+V:
UAd+6ECO0[dEXIEJLW0X(U1e8.;\:(dE;6eA,6;6=3(VWKL2<]R.T0b?/Q<T\A<&
4;<_LbORI^27+@QG3\(VLDfVOJ<UJgB/MVa+HQ+H;F^d[M[TU\D?J31EAeBP,aNF
(Z/FIKK=>4+9TYZKR&2DMG.\UJ47]5b=M^S>cAK8R6KZF4@P_3\XHA5_b9.1?e&&
C@]:3_Y+:PPVL=LD/R2UU0D8a9CW=&<#6XS>O9^OM.LITM0?BbSUP#V#MJ)J,N;H
/RIZ8UbC9HNg<MfK\BB-Q:V5+#(RD<_YYZ)K9LfP(ARV9FHB6+Xg(b_R>->DUfE.
d)V9CD,dJCQR[4[ILcQPV0X+cMM7TJ,O#_/(F)L06_-GVT=O51D#aRKI^4eD=W4G
8^cc1/_g.U3A)N3;(SH.T1CZ^W7C<(T++:SF7WNJ9\g[[PeGWFDP_Qgf4P[NgOag
G7b&E7Z\(H,d=-XFW@.&3L@LB.C6ZM_0,g>gg9Ig4\;@S#g?#3AM+aB.b?WIE:(N
>B(XE(LN@P(>6FLb&)JMEA16\;ae>/PgC+M4E/=VD]&eO7>H>/LFa7DJc#cB1G[f
..Ab8@X3\+Oe:H0D.A@FJ-5((HgIV)^LD\4#c?I^P,3[M3Wf;-N+[2eZ:[I>R7T/
X2,UOVA/J@;LDR9=1=d(0<gR&26H+)C+T1V(7-e_Q\WZSXGC0=JK_>?d(LL@2[P2
+9Wg(I)W&L]Y>4@U_,JK@,U5GXO4O2GO;;JCBI9#FcN44E[2^MdX+0>.(751B)U\
DfHWDIRIV&If_93X6Ef4cM+#8g/9[HgJ/H[A(Lb#+PWf?W6[,_Vd3,A_1?LW605;
.N@DTV=)aUW]P@?YH?=Y86KSJG<c=?HY&]<;2D[W)g5(5M<MA(0-0-JSOCY]+O<e
:J(aBBGKC:H5?&@3(aN6+.=<#]6&7#Cf,VT<5@b]720HR1EEY72JM)SdbPK.]29+
1\@]/OX\;a+HQ3IF_@Z^PgOT3LL:8[#Q[GXce95.5>F?F=W&V(>]2+W<,3+?]<b3
G89V8JYe.DR[a/a)VA^@Q.0F/=HIE&A7N4YX2Z+I.G@9=gS-P>.Q:b^.B:6W?a^T
4C8]F8W1CAQ5>/@IR):^C,RAY#E]9>Y0?OfA-#dP_UEB^QGZ(4@+^)/JN,[AJ?Tb
b[Cc=Q3RXIE?Xa(53FKANC@d[;=8g7M8JAY:KM[1OJBY;fee45@62f&8&;a./J++
I.9V-UCTTe<P]M=[]?E)[ELH]Ff[RFFA#RQLHVKV4.LGFA^AAJP5@9NNV@dG_XEF
025PQL[O&47P);_BOcXff9T#bX^PBTc(a6PD)ge=7g+>>CaO^CbE>X47WICD3QVD
MF=J.[X1M<A8---?&Q=;9YW+Lf)c,c+D4MJR#7@CQ3e=-Xa,b+N+G-aa9QKIBP>F
.WT9eAb[/Z[f/9R8-)_\99DX?M5TRWKK+-6_9O^bd@KY<R5I0-,E8H8eFbfW1;46
.T631]7/A^/J.N7TCJ33Lc\AdYQBeTJK_?B&2\d0SK/M?H=8;-bXWDdW2A9--YYX
W?Ced93?S_M<JUJ,R,:]^1f\A)a_42f;S+W-7=K)1J/6UEXA<7\eP[T&f2_ZC#G@
V.b_df?(\Qc[AC,_?<gOeN,T2+^4KW73LYFFL9T?TDb0KK.+PMR8c]WL83:YB.F3
:5&MRAN#]7gX2K,DUGLfZF9#;Q(QTFH,^FH]H^81F+^eMY=W8B00RLWS\:g3be;@
G]T1?V2KIGg[f_B88G\F\W7D9#22=CXd/JZ#STW,cUYK?2J6U3LaAN@4_eTgDQB7
3O8E1T43f6,(UZZQU_29/Z0?PQCGg,&62(K0WZa:)K-/MO>N141[?/8Cda8+(+#J
>NYCF#F-HF_Db5WQ(.TRA/Je<W7;63Kf^bY#Sb\R+B<NYB>g;)9#LJY?PQ)V1TRF
H/?c]ZeY=(O=;K+_0&;K9UZ,c>@OC,DZ/182N15P?Q=f]Q?JC@]e;5cRCRZ+M?L]
XUP=Z0,+7B8S=6\J8)D\)[9c//\,XMH<U:O_\a7@5EI;PBAEGRKN&SNH2]XOaU7@
]WB9U6.G/Z.KU0[CKL]J474A1-/G(e:477ZA8,]g=-89fKg6JI#Mb@&[E=A=&.V.
,MI\a&K@?F#a,3D;<,)NObBNQ36[&=&OLeS(IK:c)AZX[=L<G(5OVcVc?,_BFFRU
R>4dZA69W5P>cLP7,.RH3]76-0MWgMDQWOZ8,X,.ZPYgS;6H@WEeN#)&B3.O&;HA
3:/G^_RU2R?]TYXQB-_OeKBB08X_1Jf2UPgF;:Oa+D?(=.K^)C-47MLJ5=4PO\N-
R&E8-3[\K781dT3VeWW:6G?OF_EC7-R@NeX18@ePXP4If+]TN=FD8g\@84&M(OH/
CSKN\+M+5/-3;FLaV[GM69UFWfB85]Y_N::5=T_)]T=eC&LHaJ-39S?P/EH##(R1
71c:(Z6#L]fO0A\eYgSRV(A\HP48H15O:/U5JF?cF/1UX:-Zed=K);H1fe8>INQW
0c4BO;NcD65:Af.9Y=fHa;UPD^[[&gJ,[&CO(QLPQX]>9)1R_d[U1ZWB22D5dP49
aV,IZ<&P12MDacY38CF4N8GA]NLU[NZWIXR]e5.QZFLR2B3EJ_@(X^V418.RWI?-
d<:3C#HA,7/4:U)cMW.?]F\44\O5\1AKDRZW\Y(g#]3LAP8<R8<P<4d,&e6X],DE
>O:<7PB,Y:SeT;D]C9RcGfA,YB;\71_M@8Gb7MdV_T-O7N1()46U>2D;MH1aeZGd
bJ#Gf3AT(72)CRRL8NVARIab[:T\>D.L7g5d^-ZEXFZ3FC2E>f?GYMK1JO5:\.6W
(A+)A9?RQ@]B9QM&8)??>aJCb<,.P\WK(BB(TSaJ9X<2T3+T-W8U_DcSFN>Z@d4J
Q=<V2?\WLHaT4AW9RAP4f6TE@.dQGRO(05-MdJ&ABUSS;9JfVBH1,IdL1eb>O.aN
I_5@Cda+?K@Q1O4D#CURCQaU2KDY0OgfE5V6UCg<&MagBV454O)eJ>(^..a/HEKP
@2@=/4VYTaZ2AdZF493NCC/NA_FOF?f1[K6^R6DX)C_7KI1CgJ?+e;J0Ve^3EQS#
BW1BAG3e,/LV)MG-))I\Ub\@62Z,O/F-BI-J7[X-a97:;A^JR;HW_0+0dHT]QK56
a?D76WgG2OVB7C-@LC4D]-WDd1_U-OM7+g-T?[L\3W<OCY=6SNT=V>#1F>:aDWOT
c[E-+Y\,d.ELXIB>CZ^=J&/W#_?]TCE)Ka(ag]DZ<8HU^.;M#0A[ffbDU/JKD37A
8NY(/NZ+bF;U8(.d48#I/L>:ILR;)&XU8V5]f\)=)&]1(1?N604;@:0.HMF\1dNT
fUO)>9NLZ3gaM/L[)/g<(HQ67P2<[Da.=g>?g?8Nd8OG6KDd6?^Ka8594[4KU)F:
)RSEUC_.\;bQC<OJ0N6YI+[c+4#W#YDTcE.+>0)#5)c^1C>OB)+.#OS:?M.+G&4#
b/_7[<D3#M+#NAe8AaGK^A)=Z#+L2\U=BKgI(>\7X=1;V+C[#=ZVE&&J)_DPP&cP
2VRKPZ)&X&A^2GLMS:ZH2KJ+7&4KEcdb6b;F;aV8W_)Yce)d@)Q6bCEGaD5aAH?&
9G>L6PbDI1XgJ:<(=HJD6Bfb&Q]QU)=Yf4I(2/3&CSXZE?,KZC^(+f>P\T-QN+99
7RUACD/SZDK5\QYMTI[XJ?G16HZC/d)H3MH5=8V077(ZS7+A,ZTa-e>2gD#R(1fJ
6c]G-7PQ6X&7#dN+ObgFaM6)5-c:.#H<2);>SDH;9^:B3]J<2\MI^NA;JH+#>]gI
eV3,gE,94XCE9/P&=6P.G(GH^3&WVY14ALdWD3;[:0^3WZaFK6?(:[7N=?TCR]e3
?9AT#IPV\V;,8a9Ng6\aDPAUKKLOaT@=Ud#HR4(790Q0AAK([\<>;)D9M[LCe:R<
20S=e@HDJP,&]63d392cbT^NE)&9eb<<c)WG)]&FIg<@_fV;ONA]C7@T-/O5Ue]-
D&7Xf0J0MUPbN\L>aFZ3NF2R.IE#)7_[?92b.H/9DU8K#)3BaZ8^[ebPKRO7T06G
[F[]eZ)26WeMVP-RZ]HR7I.GB@Ff9G-75Z8;Y[^aIcLIP8^2M.9eJ1_Dg+4E^(cf
?S8Z@JXVSI_fKa@36<TU/@AOB&4-9=:+V]J_U<)Gd0:\L@;TEW+0KSM+]S07)d@J
,^Z42>#E4Y&F-EdS1cKGARLQaaQM9LIC?&NKP1^b\<6<=OS6#?N.NB3J[88Bb8T6
N=;A0D[A6UYV0Teb>L_NL)5fF(Q=E2FafU944C&?4HU+@9O+7HY,(_RcAX.(eY)^
cGV,O7<GK/,3-P:A4X&P0KbR5TA)Z&70eTdZA(GDL(ONIA,7IaENR-bg71^SE2.9
G0>-Y,=(U42VB(XSLb=aS^eUJ#0Q/?ecBdV&VHV19Q@2cW2YgZ3&-fS^C2RSGW5G
JY0dFf0.&b-(bYM.&d-#af5Q_H(8I\+6B=,CgGI/IN?M?8(;ISbF+-4d<L>]-+gb
CNd\>55aeRV-&(aF:AEORD<V#S#TcJWXT^:-98g7TLG8>W[LEEN,L#8?fZZEFa8c
JF6HS^#e_8TW\&6I)4C61B.Qbc=8)3?0^Y1+VLI547L8>=c/=/@AUD6\&1U]E-M)
(X#[F,W8\>1E2(<:E8X<2]BED13fTM_cD.G&OX5HI;Vf_6=U]<)N;.SL-^[H?U#<
FO;CJ@2e?#NbI#Z_O&.Gb=g/;=.X(&/Q7FU0dH,M>-A&\2>.:M_?X)1Y9N_,\D3/
YF8W8ab?O1JIC3.FFg5B1<W)[fc]NK1_7RV1D99LDU2#BUC@S#2AV<Z8G?d<b75Y
369YL]g:G@aAa+.VP:3a6,d,NR&3PGCAW23ZafFN6a04[Z^<-\OKTc<21c_b]E,D
#<L,\R[>\/\Q1VXX+0[&5W[#b_957;73F;VUK:I@B^/G^27MPdd[/E5)K/HOd7BW
<(H]?[?A.@b/>0)3K2M(RL-+bdQBU5/b9YDWVGVVS.1ERafH2\g[1T^T6cE;\.BV
&;1b->2Hd5b+7@Sb,&<]KIB-@>f&FDd7QfFVZ<\NJ_)&e3Z3K71<X^L4PcYNO6/1
#WOE#A]cULK<Q:H:,aA&8J]+)HE:6WZS54I3_0?D..AK-\:>WY=J.1@/GQPSOdUA
QYbBb.+]YgV8GVOMRQVHF,4Y(-79]=OBe1(::&e(E>(S6V9bIaD)<.9.4JG)<QWM
)>K]KYe;U6NT8;[76+FG7,IfT(;CW&+_/@dH88ad=V7Maa]eJ82=QLB<aL5D\\CL
dB:9ScW+N2CcY]MPKQVQ^A<R^c0]B4Y-YB&bI/EWPO_YA[7\WCCQG-UQUgSIMe2:
,1@VX&E1MQ@INA_0Z\.M-L]-Y3EOIC+9OWHP?E3)#.A8VXEOfO@S^2d?D+V#@(gD
5A-CFJBFL+WF2dCS[#]4d+T<5,fNT)U\.^OEGVRFXG[a)D-@a^>YPLaU_FC^DDX+
eeWN>DZ6NX98+gb4E<<>X^=M=S&)e0RALJ8b-2D;VYf?BL7dAPV8TV4;.Y]LE-41
3SQV=F-7D@;2F-[bY_E-;KIdg9D/3IBY=I+5?.bCY331,Y&Q3Ba.d^0FS28OZ_Z(
8BbN7)IO;df(J=2)\,;@U8[)6/B(\YgJQOTeV,+^D\?;Y,R)^Q0>.@HLTJ^T#E+Y
WC8OZCe(>,H7OYWZ\/d9&@GZ>bPab[7;VEO#U(T6>Jb@@Q]F:P_B-&Da[VLGf>XX
CZXa]<)QPNV0]J[J5Z@G/b3V-0/3@5&RZ#SFfK@8C(W#C?g:NB0G@M.fO23<]WCb
[4+][=,2SdC5)[A_52?Je653&A8&]#^f2HK3AOMdB?HWPW:d4A:4d#(QJX4;)G[Y
(V(Y>>,#PSXDNH6Q-d8<7>BINTY9E<OcCMV\AN5bPcH)T(8CC@H4fRS??VUE<LCA
67EP)?=_(6.B]K+&Q)#H/)M=9/_fWK9&^+S_b4,Y#]X>3N(b6f7NAWJ:Xd0X58fN
Y:8CDa)>EGO4d1?(IbfSB4/-L1e<0-gZ+6HaE1TDF2&I=(d7RS9LdK;KPL5W4-?4
/Ag,F:,QVdGg\MV@77:bA):[&gG+>f3B]AR0<9_2?g1e&D=\fY\P(L5EWEb1<YV#
3Q+H.V=<SHY0@eOd(Z[;a&BOQ-YQSB8Y:L>\V&9SHcGObX]GSN98YD?R5)LLEZNK
GV.6>J-&5_&V0-)eRZLS6U@b_.GWE?f#JP2]R+HQHQR.Q.gH9NaV=K9bT/&I<LP3
R]_aQGY5J0ZJ@(]@c-6^(#B56c.S,76RXf])_#90b#aV_Wd-I>C_<-7M@^SZ40(6
f^:1#UJGaAV+.cFVS1<P9A\+-B<IeD](DS>)Y;S,NSNGX-aZ(3eJ>^L)\IfcBYKW
RSCFT2)AE)=4+P-3H7=eX5=.#3Ydd=E?Q#;G0@8.+bJc6E=A77>(^4ZV<96EaV,V
Rf0-3N9NP8#K(d#Z\9:If6(39&F?TT1SbeBBVUf(=MG+;2G+WTJ9E/g&VJ]8LG:_
[eM>g<A5[&.U@.D4I3CH8L+0?5[_,RY)@19<<[T,^O[V=2=c5ZE2a5\69f6B/6/;
)#gfKQ/e+/DE[Pbg^22[+\,+TI<39/6XZ>JUJbMIH>N>^284>,c5PX,^?]:4CaM0
T:aKW#7S]HX857_6cf-cXCR0=YY^EFD/+E51B,aE1NJ[9&LW<cXC=Y]_,IaTDcG>
7Z_SQK1PQ8,-c\G.Z8JFH&0HUG-CA:5DfeMTe=,&a<GR..g.H,SA<fC<65O)Af,b
(Rac),D:K[17-MPg#&[XFe,(eIF;<@fWD?<4EP08N8U5W?)cUf6f(Kg4)b7W4;Z/
J^_HXRN@+1@c0(agg3We]P)^(DR#E?WR4OT?<V7f[+\F[-bOSE<S]_/d6GXZFbc1
b2G.:-,aCbL-FUE3aeG3Y91W;VK+A/@Vaag6c,[Ba4SeQ8@Pc#3;W=5_X7(=TBed
OGJ[Ab1]5<7LY/>^5OMD:N;a5AO@fb1..:Ae\dXHgO?]LA/?YVK\JPMEY<6M9:7C
ZYX8_3^CL-c1<G1fO:(SD;P>U<V;XYC-^^\NZcdg(C/N#[VL0(-&&=0=XTd9UQIf
UAWXUJ;.,-0D&O>YW;TMR.6TXd&I[]S0f5Cf5b3LA70Q<U2NPSY81Q1E<Ld.eE/O
T,_gLB)3(.Z_GV9G53;5M9-^+;/?3=F/SSS8XNb8VQ@cIK)LDC?;Jagg)@g5&]C6
\8GaS-Gc.;\MLI^V2_QEPXDIE[H#&]L,,\?^d2B(gO8MJP>Ca)(;Udc<N0d1(Y?4
F4Waa+ASAP/0\T8SeRVCVG>7bf#LaT&Y]X-586]YO[\>2DeOE)(9\JKO5LO[IO9/
F?R)We7\:?P6-FdYN?fTNF:gX_b3=D@<7eA4@CT@.eP.))[FZf-<:/3H0B-+>TGG
/00WNd0?_H[Y;G,SRKA]SF>fgQ#+_4S73aeYPT/;U^Td#7?OZLc4\SP]:dNXH(J@
TBJM0BFdM.8<afM=\L^g:LCWfM=7O;KGc:QfDT1cb\gd_EW7a.cVgD.8;U-U^VB6
H+>(M09Yg\K3SZ,caQU:&O29PJ61),<[\J3J/2b)?)c]I4cNVI-R&gVJ2/J:0-&S
7PZa.31C,\5>/<dd(DH1IG\5de4[ED2dFd41/e^KX/OCBW_(3cZQRWeWeL;0Q<<g
>,&;VT.[-=.S4(eSJ4Dc_.M3LPJ&-\A57I[J[c7G-76f_)QSNJ<YL<=28ZO2>\0N
/2A]bW(fIPbY18;gT-0Ha6c<[.]/+[OS.FI9db#A]-<_d-1PO[.T-b-<00;W&(RH
FC>7Cd#+FH0OA2OXN4X<]YQ9RI2M&<&QE51,#eBAPF5bUEUdDabN6d4bd6>7QaIg
/=LEM.GD:+VPT+Ha=9064)V@[9<CF)(&&Q>2PLH+^GO;3QZcFS&SNI8+OVTQUT,:
,Pd+C].)_^gTBag6M,^+ACR)]bgf>E<SEY1DDS8e8)4(^WTea3N1V4E^L>EL<1)W
c6W1?H=<@33O;b,X>8PE);B3c,J8@0<)c@C63DN/DQNDE<7JeKJaE5M6WcbNWF6N
NWX8(,BG17N(&0de#gG_9@6[ef.V?DR7\),;@f3;ZGBL?DVUL[F@P>#6:aK.U9HJ
66IeLE75##eNSUcX-IM&KCc?WQS,HO)GD;G=aIf,H9NC>(ZV0WYN@Be03Dc]]VKO
1T@M^b1:)6IZ(A#ED[N1Q,76?#@[c;DIaBEQV93E#D<F[6g#ccC:fg?f4c9V7#+Z
YJ=&)>U.;<bH87C#ecL[0IDcB34R\J43A=b,K9Y(KWJ1M8.=&-46Yd^DNE2\(f^F
_1]_fX;I>9(,f+U1QYV&&8#/TdIQb6\H.7M0JW,IH/?<3Wf(JF5])AG.b9QN_.Dc
d(eTT9,[eeKT1ZI.W/T+1&?:Z[2P:eXMfOKP92/LI.BL^5HNT=fJG)T5XFN.Z3E>
U0Q.fG@6T/\>5d:DV^TE)dD7L>O()BVHFWUQ);;#eLG5]?#P<)>cJ^:\&@8GG4+B
A6E-><#[2LK.,Q49>+Y62CaLc-F,O_F9HNaPN^@3CMg;C9-Z<ESe8,@C8=I#649e
_Ufc)J&.#&A)+^dVXTeNL+d/g\JC6)6bHIX4O)3F/b]dFcA-U7,@70O+2S0.#FcE
cZD+4ZML9/_aQ;E.HI=&])fH4]7;FCW0f(H\IES+\BI[DHbAR=[Je:L^^)N](H,-
@f.=,?O^),#?#,:@DKDJ:>VMS)e995Nb;0a9AZ3)\>08:ffKBGE<=d&3cD,Bc5-5
L(ggfBO7D0BX/6SOR@PVU>^UQI>Xb9X<?\T]^2B?GLEbZ,?],^S<WZL>/2-G1O>4
fg-=?K^BeAHZbH3FR-^WD/=,MED;-B5/?b5[\OH#eNOXNNeL^Qc_]:FNFCZ=6d.K
Cg.ffHE>ZY+bI0=g-HI,(?Kb/dAf7A=6K._ACW/bG+=cL-)8#C1E-6f,B/#<1fg3
G?4-)3KIGFZH5,Sb3b[d^AV26RHH\f0>E-4(:^F<;P?=9E]/UEUdI8@B5?,\F].0
\T38.NB7e#IAY3KO.eJcE7.8SeV<4;VYR4\/CK0=+)74AL.5fH]U6LVC09X/(c&.
SIRDPCMP@71La4P/Z_7YE\9fa56R1S4/a8ICNB8c=T3C[(a^a<5M@Ib.N0SWPfL8
^DJJ0R]C:K80-(c8OP90UNH7c?G<)3Ba#3F<&a[@OH(T[De(-A^ec@9#6V;A0e^^
I8@5IM6CO-/-8.:75[GNQ4@=497Z^R<>U)fU9>KX.9VWMdgFHOKADE^)1#gGN,KI
(QHW2O1ZW0X>a<TBSBEF[e<0f1=_TRZgbgEdO6S]Ad55J1SEUbP8-E55(^ZF7DKg
TKHLgYF0ZW]1],;JGCH@XAR-VLGYC:UO9]4cM2@S;#V.3@1PBc1ORd+GZJ,)W#<=
ZFY,UC3Sag9D.OfLFdGaO?DMQLb+_^2/F+_4<[]@AOI^VFd#cYfK1.Ze9#<.=XXE
X+KDG)aXQE=[8#gW:b.@Bf9/I=D_Q+X\Te6^?5=FBOKOYad+O](>N]?D>PE#F&B1
S><IL_42-[)H)^W:K&HE-32@[,U4I(.XSJeTF1SgT1&=XQ-Pe.ccRF^cY\5P:+[9
ZGZ9WI)TZE;2bcR-FIK3ID4CH-YKc+BVIgY_Ib>JD<-5/A(gIe9WAYVZBUaQD?a?
A;\SG@R+:9e31@5X^EV:d]=2Y>)F5=YK/4]J8XFW.USTEDSS:cI>Q1.->-01S;(B
5aQaW#BS]B?C\[I_)6=XLT6X-P40U+4aOYaeZF);,2f,F=>TNKLNeMA(M[1#&32L
2=0U+K5=^EHV_NO9?3)K+)fWddNV3_;(4K5b1E79_;M4=aJ4,eBI&+A&eF5ZA18B
GF))A\LGMNJdd;U4MX:0eTSLO)5U3J+KDKHQcWPCO@^7.5.D+3M).155\B0XKa^^
3gSf8-ad0(C(8e?Mc<]D/J;-_Af9KT58(YWZ2U#K]?1I1LcJd-@-:ag1BO/,Q^[-
^IB4RXV86&Jb=d.,f<_4Y1:20#T/VA]P=S[^B^4>_NcQFNI;-@_V,fA7g^RVINNU
Ig(H5ZgCT4&f[1LW]@<b)UGOC^@^>28,N9B<g>49LN>-?Ec(/WDNQP(:=<=&>)I6
VeAX#B:a\EECWTA:WUAS_<HY4B[_GWXVU4/^aC-<[A3a7_1]1E65FACZ6A(-T/bT
0,F7G[+KEf^WGGD7CYgQJS;ee2((7cKU7T65TT?c9Tgb6^?]NBR@DY5:@<K:>H[N
K:L(\(ZD)2)-J;/\c,,fb._MT:aC[GLL;71&?T\62+U?9&E;S,5D?0_0KACTeb<B
<#;N;NL2YU>.Y6<8e<WQ]2:>#N[Z@-,7E:&EC8/N;=d(>-M,@>Y[Fa./eD2<WNd_
;&WM+UL4\?X)@3M8eKW^7S]Z=4ga1K]<^BAL1SR5MU5YSBfeCN[=:GP)e9F8e4S2
34E#fOS@SB^?8FA7J1b)+WB2--FaI#G]TFXEb5d;8F9NAgB^3Sd1INeHW=+CQ56,
?aN]U:RX0aA@L0+@L;;DLH09K#+7:U&eeGI)GeJ3=W2)/^?XV^].W)f:@^&aZ1+c
;EdMd/F9:7eE+Ea]2C<2JEJS0P9eKO0(99-?<O9#A&;7X9F>-^E4^H9M)U@_?#;9
-M<+PA:8AUCE/0J&gE>ZRD.IB,X<b738)M&>SUS0=<D?/J+eb/4)SdO_1_2E\.<c
fYI@4<9Wdf^]2>I]#AX=/1A,YAN1P7g]dH>(+M&M&d6<gg52IM6BM:L,R@I@SW_Y
2VC,e&8C(H<=JXg-.]BDY,fN8WLR25S=cZ;EJIO;Wa6Z7+K[ZW6e9CK?:L/],\a5
-EI#ZbPS9-35S<(d@,0TeA1)I(V82;T.,^L\C1YM5(fc1,5PB3Ia&UW9T;4-4]QV
OEgYET)R[bH<8\L3<>F:?cg;6<MPCDfcLB=8RU&CRC/dN]7KO(2Pg/Kb-:2c<+)Z
IGUE.X0gc0^GUMf^\fbT0J&&ZI2Z[F-cTc0\9cZC+_f8C7QVUW?e2<P1#cW;Z@/W
gC^.?1;]0.#KePS66\)-BBYGHWOf\S,-)JF:NMW.ZZTZb;H_6GN(RO[0^CD9c);+
W(g>J,BdP>XNdWY1\Q9g-6R8[_)c13B(HL2N/+d8B<g<K;HGH>^AC&Q:03dg060V
<TWY<A7(;@WXK8<P178DM13D.Q1.E5,3CZ\GbL=._W,>7K+F4GX)2d)9S;:ZcEI,
.gO9-EKc1M^#eb_?L1KJI3I(/DJ8I4X[\ceH)J^G>=/E\+;ac<.Yb/_P?N?LP1=K
FWZH]/2/8KV#?R]U3^3+HV2KaZ7P]]W.e8UU;M,]9?f2=aQE,J]bW(T?<K8N?#[K
M:3G=^&7>=X7LTYNHKN?Q(a==_P=6fU1b9FTWUg:VRIQ/V9AKJOaYQA@#=P+_]2A
<Qb)8K+.Xd0YA@=5:PZ)b4,H=98,d1<FaRS#_f21.B-I<MZbe(WM6<9_K:^JTMH6
^HO<VRPN^Z>J0YZ@\3YFIMCZFFYab8[,(a<707A<J6I6?UOMPTY[L\06NgSYD4-:
d@6,,UY)Le6VNFB]\T5ea6;@1^,4:GA_:[NG7F4>R\fW:aDO&g,OBKFA=_JD8SEN
=>_#(KT/.;2A_9_,0C1\#91DFACN5WZA#eC6V\ORQd(A5(a]](THRFg;8QF1LL<F
VggOdaU^B2RdEc8=42\]=FLQ4O[W_UO105C7cZ7+Ub]M,#2<#6?B-4<RVZa[E5(.
Q6/BdTNB0J3^g80M+GcWF#)aWa,7d(1Xd.((HK5JD[\1/5@T&.7c7J[g]33=@WKL
@W8J(/EGNA4I(d>/#<XZ99EdWBOXW1KTRLc5]WID#Wd5?KC_R69.VD@ceLGAXC/[
+J.dE7,a\G-FaLU?,4_H30;Be^bJ51/(db]YKBbY)daUM-ADSK.[PgDK7PK/;dZc
HW)c[5L6P#3AQ<a#ZY,+@Y_-.?WGWdCX7W>EQ_,B5Q+,&&LY1d&ZG4Geaa<5gC3M
S?\f5bO?Z,RF0GJE@_N@5JZDGf7X505<KB+N_:IT12<?]H/.\VZWY6ER-@#=[Pd)
#[A.AR>]])K[Q\,R)+/1FN+X\M2S=3];g5C@=\TYg8FDa+Z.UU4DXIVZ3?,P:I;E
/F>K<]L-L9-<50T_)1&J[+E8[&g\GO\f^?g/\gQX[[DN]IbJ1XGU&LB3]GY=^K-J
[(+:NG>d#R&XX<8TH-<[L>6E/FT#,YR@EN4TG_IDL0.0VH9P>(Z0<6D(VJZY[b,f
9e&8I4@dDdH7:)6QBRd9;;=-3Hg)]:>D6?fLQ#TL/+-[4/7::V-g1^G0G/T7]:SM
MAK=e@LMN&:/>Ga7e-#cDRD8A@I=@8I>af@</D4bT(bRRN?aG38_Pf0D(eJcG,RC
DK_\K:-g]1DM49=I#B#K_Zf?[4;AgS]&6gB8N3)1_=__PWbeeD#PEVR,/.TDRK++
g@eYV-8O8VC>4LD6(A/VFd5[@P-c=BP]O4I2KV0-1:KNE9TQG_U95SMNgB)-BIP/
:BTXIeE(6C@MQ7(G1e<Q-LAOf?TVf^P9_KW\YObU9.R8_G4_XCC\c4S7a6SDVR4\
S>Ya5_E]#DF+Ba:G[1#dI@/<D0324eKWLM=1ccC,+S4bA;gZNA]21Z\CSH8_2F&.
&0P<\B>)57]#b.U4+S\K(Q.Z<3P7d@3/T6)#\\R58G8Y#GF031TUEC+_.6CJJ;E#
BR#F(L&.PN19DT;=TEL2@dS9E>-Q>H8[CMGJD#FGY/;V[B=fH)T<c[T&CQR/<720
K:Fc,&.f5V-?b8@Z4GWS&MO74@,[+RMXdGZSWVQP#PQ=[1:0AY2aG,&&4gG6:8<.
1eM;/8X9#O]E<@._?,_&31=8XV>)FKK,8(]8J8d,6f=^DbICN2M-GLTdVY#\/;A_
-P-B_Y(2c(b]4SB=1;KXC46P1f0.(0;V\C21UA[U,Nb??[(:f:IR4X/D0UPL^\_K
-;I;01AeT=f,1a6?#;:T:U,Fgf+Pe>e<W.W)5]M[PVB-Cg(MK6CF_5T4E01X8T/d
^B103&.)Y<5:VcQU)[6gPOMg<:_FU<6KA0N#Q)g-;R<[9,LG>ZJ>Z(VZI7AQgS]+
d7F;UOaL;ZU-ZH_?;S(a4:H&#e;5KcEgPbfg;(,HbO?,)G:+b56NRMUaS?<+YQOR
0C(F-aC4+e2I9fQ?4I7BTN6N[b\=NTT+aMOO:JA=)_F7G#J.^S4P^N?0VMad_-g/
9@eNfH&_gKW13&C,7Z[Q59+#@TA.@K<D[QbT1]1B4JG?T.,C&][Pb4ZUdT(R((Rg
DW.1GNfC?(=HX#b,YW6Q:M/?4a24;AL2I4T+Y[.U3<^[VTcB,=Q9bZK9WcX7RM)V
=S:,&QaUBP1EfB=8(9^L(350\-&J),S0b1aV)EQ(</4]:(T^[PVER<,)Q@M<e1c(
Z=0=D&OQ69(7RIFWb7VPVR;/P9^M^MBGIL)@=G=P0F6_@K/7I5AIU<ARB&Ie+Ha;
,5YYUZ,U2Zgg<##BP-FVC>:0QTJ6SJ@RV=8.0.[>gH0L@8.XScI]IN\=5A:<fV@=
?XQ&)Yf9B)5K5:b364BFE#64UX1:/R7G_C2Ge6F?eQWY^NF](HR-&]3CG8&:P<^2
ULPA7Qe=LY+6Y6.^aC-B+Y\\9,YbWbaK[O4XJXGe)ccA<;^D4:9edZV[;UV1,c5;
?_eS]^K&#-85-0Mf52J]:BN:\F5KEA0Q&=1,eGCM1C?cH&S&S_398JPI^TYMX1.Z
-SPKN,?P0+)bL54V6RBZf&\DEg:#OJP22f((aA]L)[Q8W-FA(fLZBO8B_#_e-\]G
XDc(J1<&Ua?D/S9HKUf;OD^:#>H8L\PB1]L3>C96O/,99d=PGe5(S>X&ELM(VQJU
>XG^4(2:WZbL4+Cbfa].VN1L+D_&T:/#M[P>N(aCGT@BeJ;C_N9-I,Sg[.d?.L1M
=7&cI;;\0H:>R^A5+]A4F>FFa0M(:9VCEbcI>64g7Q+F@NDe5b1FA2&EG9HBeHU0
X2T?E9+cZC&,P@N5=R79GWV8;RCHINX[O4L&G?QdYeb7WVCJ=^Gb;)fEZ]CK)WBG
NdA#[F@-UgAP7+<=&&]bHV:<S5fgF648R#g>Z5.BAM;.>Z7&57HF)M56GJ\.g0e=
Q(U(,2/J+bJRC(CdK)eFc3NUMf&)?I0Rc:ISaU1Z4ZU:J(VI:M>V1J<7H/Gg[F^M
:bddOU_92=&:a4NE,,O5C;U@SMd-?;]>&3S\Ob9bUfAfYH04Q0BRUdG<]cYN7;A)
#(W#R_K..KT6R??(+PE6UZdQ8-7H8fQ4Vd>dAF6FDg/>L]#[033UTOS0\T.0[4FX
Ja<c^4KF#J@/edUOJ?6QEB9aI/D<U<SIPL@[<8IgP8NK^aSE#=KD,(U;)BZBe@I>
_VaWDU.+JZK36baYgcQ?E8Nb+IVAXM7WbLC-g#MGQ[Z2^\fO(5D2,8d3Z6ZIO53(
3&\W:dfD=g+_H?R8KS@A/&cU8)?1/SD?dXe(JW<G^IL,C98W/<gIU12A\-e;BEQQ
\4^(QIXA8?bEEK=JdEeR@\QWQ&<HbEN88Xb5:N<#0.1OV?BD9MVR@Gd+84Q[<&<#
&07&-8f=F^_T2Fg\QQa]\WZKbQ^aR#ARaCF24)X9K.0WAeU6(7g)I_?OF[=C2I-B
6EbZFEM#HARfQYWQ?1,O#^KcDD-NP98E>B-D?&J)=G@a8ABHMJXD31g+_2VAR_a?
UdTP+2bXBd(^_)>5UY<a/edJL7NKM5>S8(78CT\ORLMTZdA:RRH;<IBO[5HfW@1P
DF1O].a=BW+aW9/GGE?0@UdbTOA@.>R-ZP#V@[caG&_Ad/03?,0eKDM0XB7]W^@Y
I,00[4R88B-T9Q)&8ZdT=V;.D/NO]VQ:7=Je-X8B8g+L_U31);;,5+R.U]MZFIEB
NLYKY27Z(V4fR=G[:?,2,__UHYJ:^,I(-?3S#\&b-+/N[N7a1F,9YF].,\O@X^0V
;DSdHX@C\>eNeW/D+]9:^/O55H<;AT?.4/J9<C:+<\8-5WFdV8AK8,<b@7[eW&;A
:B\gX7UeZ,G=2gAAU-FP4a1UZWGU&,^)<?6).B3OY3DTU>=[=H(HId):PffgL9?]
&^Uc2a:2e>A9M2A;)<GZ:G,?Q/6\6;X7NDC?/.P))/[(-<:O^JBbZTW>MP?ATH9b
aT-F&e;7=&C40U<6Y;<NfRU)GIW95NKLA6?FKJ#1(<.<W+4UNeEb7DI(E<Q/#^2M
((,a7Td)beHX)Ga/ACJa.e&O;_QB+.;DE?=G/Y[2e]KUP>98G&<-[IfS(4cLAIZ@
K24gZA-X\41^?3Ue02?.E>J,C:B[MHT<LU9WWcLEAZ\?cZH/AYfBM6/D_WH]J84I
X8EKJfOMS\NZNX@S,47&T?Y_E4P,QTDf+:TC.&R-4MA6=0T-e6c+d47>AOK<IL\E
YA/^HT.0dd-VA.K#W.PH7g),LL[38+Pe/Geg]ILa&<;C+ZX<.(TN+M??gW]L,UI.
:bPE&]fK>9PZKSC-7((1Q6,#aEfQE3dJHQ@^KV)ACI1RZf@Z9.BVc_EE00gg\f--
J([4K1SHd]<5LO/U2OV/@<>UNQ=eV\F.cgTBV,M)-KU<GGI<]b\,SI^0O,HCce;+
A.FZgdeH5^H;G@eP_V3TYP/3bcaGO&=6NN[^B;:83K?^.X6JM+T13/bX[]3[(H]C
#_-XVMC0>DbQ_bYaGg3O;==S_^\/2;C;WK7@>Z([;4V6^I3=6f8J:+1N4fgS5/0=
f8D/8IR\Uf3CMfJ)Yb-<E3)^7N-1(078<#O2f)YcK&\c4&d[VZ69[a7Kb(1W(5dd
.[YSZA6\T4P]C6H8@DIP;EAS2caC5P.T&0W4J+=EDYZ7YESYXX=UNQg-g>459[/F
,NQKeGAIa6;;GPTU:EJ)=+JL)F)FGE+5=e;VMQ/PFeK2Yc4P3Y,I?YaZRcCI6TKF
(X\V@81=_g4_<;(a@1:5#^8C8X^@S^e;R+(X5&.R5()eFg[N(0+S04)(M=U&6VZJ
C1RT/0?MV8LeUE+8HG50c\2.,R#Vd>(+7f\64:dGRDb#>BYBb0C)Xea]M[P23Z9)
Q0O<T@6)RCYK1>HO4J5(J1QfPeB6;Zdaf58<W&)^.8BFSHLH^V<eW5<,4RA^DfA1
K^>&Rg_;\O3.+g[.CXU^6O.VX39](S#MI>WdU<AV(<Z0:bCTT?I/dG@0]V(EBJ>?
6BXf4#(<;8W?0>M+FRB(b-+<KIQ+(d_UD-68b>W?XBSccc_<7,T?N[>dQ]E_XaS\
MZ;4)FUcJdSe^<UI86D^5IPP7&6W/c347:NS06b))P;^YW4.)L9.;VV;;4f/=>F6
6LKNIIJ>bZ6)f3.GN[)7:KPC(N1=>ZTcfJ?0J;BD;NDM259\SLM8F[9M?KL#[]Sa
E^HR<N3MJdS5,AE4)L(/6X-2\1#R^D.:+?eeI=3&&\\:+ea06R_VbP=6TOS:3C?]
g3VEP7R^,QK36D4g0JUG3d,.;gH?FLab&OK]PV1@RZ^]SVUUZfMH6+N:2?H-IK>d
dP[0YGIQ^LLKK/6M:BZJF1A-dTGQX8E/+Q;R2EW#K57ccOd)FRSPE0d<\>]FfO#^
NZ]@KE^@@FJgC];2]\#RW[R@O8dT)>&g_)YS:7U+Z\B01]SC5SQ1[=SPJD9g<W@]
^6A0?^&D_4A2Z6S#fP6:E+PO./-JB-fG;7);AB5.eU>[-CUKCYQ]/XAFOU[&,J0)
5&43b^7AEI)6/EZLAOgX>Ta048TM-;35bT+IA)Q0)a[IfG7e:dT&7#CS?9K=2&Ze
^78)5ed5-,(NQfC,_0]1/:AGOB@;YAB=BeK0R+=:.+4B:\W>e0c<ETU0H=#/^K,=
_OLd7KND(9SCAQ@U>5U-2DSBe9DXDB2?]0dEd]<6f\9/IR_aSV^f7W2RJ>6GSHS3
(SZHR#EDf\c.KE52^J=SR-U5SZ35C7Cgbf6>ER1>2:K<30(OHQ;?bD[O=Jb)_UdK
\;AKYNPZ#]#<C[f&)[;WYLK^e(+U>WW7-U(Y4CS-Fbc;AaBCZPXU^@b>+UFA,JF7
@U^&)^g(<^BQ(S:g(a^+,4^[R2cR+D<T;18-=QI)>g/_?ZJ\OW1P=d[F,@M3TV/Q
K&E4>>bGG4fV43RDa1SH2&V8e9\Jbg-/L^XSJf;#\BYZc(Lc]cYD0.4HdFDAfUeH
Q_/gVE2GF5Y8N^e?)F:S>DJU0OaX]W-I#ZYG&/;1Rc4+J>@49?bM@bGM/C:&gSN/
ADMGLad56NM3a/?b<W>Z25gU@895?A<DX5P1@17e?#QN3#^Y)dQEX@AZc3g=FWL0
g:T=M/^Ab9?c?PYA+GZ2WDS3;I]4+A/DAc=aLa:\WD].>CBLUM-2K]f8@g.J:N?W
A5Z03U-e@AN::].EU59_[+,3M=(&E;I;5-?YB(DS7YZL4e+W[WaYP2U(D4_C7J=X
BSeaXe,7Oec_O#&C+b[-<R4S^,4ODG6UH8V87HgZcOOGX)EgaQFa<#9J4cY#ES&I
=&e=@[17&_b>]5AQ-bgCGXFaN.3W1Qg^^X-bFIX;J(#>ca>YSeI(<T:;b@1NSN2/
GHZc,2G:+WJ77B1]SFZ[EaP?W>E@c@;FO9=ggcVJ:38(Z6c(aZM<K>9ZAODJ9eg[
0,1d?Z>]172STDU9QV1#0RTNZ[C(WO6OP/B9+OQEa36d8C5W5NgA&/ZGVLb1B<6/
#3UA-4J15Rd&J^2<,]BNKX@HS4>>.)[T[ZeMGJ4EY4J>7QCc3g/1BYcD0V1D+c/C
^OK+#&Sd)dE#)963J<J^UdFZ,Ec\I+bTS)J<5]]Q]TYJc9J2@3@b4OC;RCKFWSNF
BMRAN,E8EE2W>P\C<A.WEVB1YC\LUE0+UJA900P+P[aVG76JIEfF.J[S/W10P:SG
7M6A8;aO23O2e@VfaR9:>C@L+\b0.^)N\)X?MD2L/4(BbeD;bMOD^S3_&:8=5dVU
A&YK1?f;B2d6^2Q[72)9X:A>b/JO=Y[+\(_J4URG/@dZeQWI,M9,5I;QRFH?+17Y
>-)]:&3M)HJ00,<GU)=4&8_AgPcA.M6BN8HY_C)K;<fM-9-8>#&K7600;PB^JM9Y
:eSE.]4@TA8bM=H&ZK-VAIF##^YGRFAgb186c8SX@QF5C)C:,[)cNb0UXg9Ra;YN
/=a.5S>DIA7]]eF>IID9FKMX:3dTEHe;?T0O]HLFR.&.&_N=C&g62)^Kd2(M,<G[
6ER]8CYFA4Z2J)-Z(5LZABW1)Y,ga7LO9J-Y[4/:E/[M0@],&U^T1fCBb)]C&8MQ
.JL@#QSP-LW(ObN39TDd,?6[CY_=6X^TJFC.eQN48@IgU/<\)Jd(5,_HER)7UJQ9
\ab=XBA=K1YNUVVTM6NVLH62F::CW:Kfb[cD0f/#?O2G?=f].HOT7P3_P[+>I.RK
R;;S]aC?X@@W#N-3DMeF#eO=4C7TYZ&;M+:>S#LD/E1BH:X=GKc_M;=V,RC0\/UN
GbZ7TcO90DFg8Z\5:2e4AGR=)W4a8Q.C/_aR=DADCSUUZLQO_AIACH_U<fHK,_5V
&KC=d6A4SJ5FCI;NUQB^I8=+6.eNBVQNd,K->?@beO>G-]X06<D6T;DF@ZLad<DV
0:((8gD/9.FIZA9Ng4O/2Y>J]JZF<D.N#QJ3_R98^]fL9KW56.#AE4<N0geMfa8c
bS_>\)+eg<cFEaP_>EUNZER.:Za2UJ9V+G:R]3g5ZK58Bd0OCa=RO]D0;E6g#ZPJ
g]8EG//_@HG-ge=<8X(I<11IE2#)).>@]/BEaZ[X8P>)FRS;,&HbQ6\2E&JS;[.^
]:aE:H9U99S74^639g<f(-.[6KW.>X,-8W(B.B-X=:F#ZKW]G-.C23e4)^65K1A1
NYH^GC#PF9N]@Q06.KZ/-=15<c<,A8f]+YW_7-87.AJcY[G:C/T[)-CVEGSFCP8K
^5Cg,)X(A2H5UYBG<13KBd>(KMS02edVeKD&DSML\_&U8)5deB5;G&P+V<9:XL#:
XDF/A?=<;L1a)N;fE)J,H9bHH>,c(>8^aOS4+[=>KRB\X21\GR7]8/2b#NM_@6.Q
5:,d>bG3:QEQQ.9BOdQ&;8X=3G>,f?,)V2+>QNd^g?c4f=(ZOD3dL]T&??CNgF[)
.#;cUb>dIGL-7_>:Q0aSOWY0U+RHJKM.H^\fY^J5F^(2@QV,b\JU?B,O)B13F9e3
Z>:;Q&4GL[,JWadZ/MK8-J,S6)X3a+=@4,VD@b@c6K]Z;X[@=M_S)cO/RP&2U5KD
LJSG)[dg9Rd,+PKH=E5K(Y(eHX4_@@aU->8>_AX-T&1Kc.P<TcJ#Sg:X<DTb_H:&
L;=f2CXQ5755M4;U:&6<M=:K5_L(P?UXf,,cQY1a\L01>RdH&I^J@ecS_d06N58A
>c8C1;d^4PHZS(OIFc#A=?IT0+Fa;&XWZXS0YQa?6E8BF334#0ee_09G9e4E^2^I
03[^\ZeB[-eM6ZF[Q,_M^>^0YSX[;=>_DcVBB@<V+>.:K5:U;/Ub<10e7eKB]#Vb
+@QFe-4:.[)N\U7c.FFAKCc1=,3>8ObM,NEC0#+\0,TP=_UIJ5T5ba+XbG[Qf\ER
@E;dO1TMGH(-<&P9E_+gV?C[2MQ,KX5>TUXN2N7Gf3cM)>K/L&GWO54/_MTcQA<L
@KZO&<+K]:F1RaY[BE2a=BT0+A,TL=^=G7dNXESLbI>6G92;76Jc(@)7L^2OGH[H
A+FKE/MM2?0/,HF(0;;c]]\H\5YROYB2WVKK)/9.8_/B4FaL#30H2>DVJ8G>MB_>
09.F-D_Y3VW3UcDY9+bA?g7-Z9NcL74RcP5(8_:;_VLg,OQEMaVX>c)@_a_#VW@7
:fR-P)Za9;]=>Q5K&aMIO8C-6g62QOB1K@PU>HH_<d-BYdZ?++)Wg-82?6,/TKK,
XIMgPI>?B)-B\@]F8V@8^#f=0P[_\V]/X<+TZG9Ca>;a_]ZWgE.?/OLgM^L-N#ff
C)-[\c>>F8E33V_#cc0AQS,CO^bC<CX,-R.(;Ba),Ub?N#UHg2c@=gEL28?,<+B[
TGD^e8Jb3DW^\)d.P&f=4XF4;9P-#@KL]#RM8UT5?+H;#]EaE:Y19e)Y0:JZ03U5
=.6UIG0>C>:_7_;[e(0&#g?:S&1]-9@3[B-K:R+gTDZ&]+U7N9?);L#SYEgC>4IJ
CEGSE(GJSSM,C75NAXJIL;-NL66:/XaDbB;X)eDR_+b=4&S73NJ5)-42D>>>/138
SM6V563\J4D8YIAdggYR^&]&XaQ@VG3B1P7SYRWNf37OE97ga>>1^9f;AIIUb/:I
GPAg38N&6#A^#;K>Y.&-9OW+E[ZC^CMB_4c3+)&c0V-^b<Y4VYbNM2&f&f9>Ed7=
fM6.9&aaHg;)_dF?AVG#9&?CaQb3QZ<5OE,KZF.(Ig7O=]26P[ga;Y?>J^+8X<6/
D+5f5(/YX_f,dD7FENPQd5<TeH5=-g?:54,ND#-OY+_aFL&Ec:KG][?fNa\UM4T6
_1\\=X+Rf;e8UB4I(TH/57>V7-QP4./JZB09S#B5Q:\)&[)A/.SHRIbN=cC4=[-B
HT,L2F9Ab?,J29:/9^,7gCI@DEHU?,>dZ(-2AfZ+0-59UGA56cZ:44Oac^8YQ):I
-YDM4BU(a[&24gbIQV1S+1NS;^)dN<_7S8Rf#/(]E6\M(b9fc^\:f+bdPE+=\<KN
3-SY,)9_RO4C5/,P8eaT02QAdeL_^SX-::f7b7;UQ7F<F8?POHcJG]93(QY?\)O0
1G?T]-M.eXV0)gIc3]dcI=,;N)Tc:TIJ?94][f2fBWJX6aLNAO=.cV7B8bN8;4Ic
AYeHS1-eN7(,(cU3&JT&gSeJB4>,=Xd^gD+1<2X(&^/9U:TMNeZQMH4OK@Lb4FeW
a=NVU4Ogc(-(VQa2QC_e9VQRJ^B7AOYI5(A1VIYXVU=Og1AM3fb4]gdTJVZBPPX2
[e<&]L-AH]J80R53e_R7WV,1?L&&7c(-Z?N)),bFD1>g3#6QM@J+58K&;U-_V86#
&/YD\c0J&RdCNbK35GP7#+:9EUNHPCXVSI9Tfa46)=77OcVHaYfD6.G&#[CTZ,O/
JQTONY?bE@JT\F]86F_0&Ade2&A?d>3dAT]eEU^KPXaFM6,JHE#)?>e=34TP1Ug[
eI][g?d(d^>\4cJ;=.;T9]:XVT-f28ZUNK?,f\aB.EN2O&A9I(4U1:CfTNHIaFe,
7GJ^F+^X376d=S^Fe;8+L<:T(B=P&-?19f5[aSdY>8]dWXETNd]@?;XL1ZSRF>@=
.[4\49[.fKH:<VVMFaf/AN^fY&,DMQJ<N(_4/FO693L>ZZ<:PMS&6&?R]064NdF\
C[NX><BLe35^;0I-2[8DP(LJ<)P(VdbH,ZS+9HD5c,L#Q6G\W^63eTW;5]f;V-Y9
Cd)K-C&&d2<,OBSJG>[-9JO([D@IH9J)Tde+LP)[_YLS]]D,>\32RDAD9:cJT;S8
KARP1F-9G;fg^(D/RAD6L32;\TNON2P4D-K5]e85[2bVA@e48;BY_KP>Q?44=6f,
#T33,0,F.]@OLf031WORa#TWQA)0M#5aVF1L;GH#<Q<d=T]6Q0\J>-=g/5H2,F(2
>XRKRH2MFXB9F/VDJH(IeR&<J[2GN[N&7P.M].(G)VOHUGXPRT&AQ_1@R]F,R,2b
a\IHd]0dQ-_/U7^@dI4c@#3K1WBNH))4(a?RB7LFg]ACe;c,;\PWE2fBgAHeSB]4
AG3TF(@0V_SA#6RTbX-.WRP:8RRSA\YX:=30]9-RL(V;5A#d:-=/YHM&HMNS>C-/
^P0@\+(0<aGBW-P-&)LgJB1;5L>-(Q12,Lg#O(M,4,?b:Wc+AbCVP6g:YTFFY;GV
?:M.(RQKScY)IX#=?3cMgANaH7((PTL^Q2)8HGb-P//UWAM7/6\Z<F-).GN_Y8NT
N&#fNU)J+0G-^2)^T^b-@4dJJ>\)+?9I2I99>&((;KKG@;;Q)4NDAT@V+)^[5Lc2
MY7E<0c^/V.a@SZGTC\EW<SLJZBX^R6=eGF/&A+K7&,V(A:g6bdb&UI^;Z/+HT\,
51c5[HEJ1=7Y)S?Y?#S21Zd([@>R(/H/@5G&:-DVW<82(DV:<LAIXFCQ5KQ6KP>Z
ON<-,-IK<?e),\@b^YNNFY:KU=_)-fg+a\>+=<?;.]5W)>4Be#3O8&WP6H-/21JU
Tb>AC.Z1b+^L/UU25N<G>^&^R]@O=[=]^XS7B.&,6699?@9d(&XLWD=7e411.<N>
FM@?/g;T](@>OM0X:SABUN2F4RSC5.;_K5^1\b^?Y6^[[[NF0WGe&]@<I)(2D[94
4-dEEWDP//_K/TUGf#DMcYgCL)Q_>Oee#1K888?AE59Q;^PO:O\9V[UY,?1=:JW7
U.U&.RSe.ge-=GEB]+[MDC(IHTR_P3Q<c4Z0W@H27>M41dC(7fZ5^_5,C,/c9JA3
Z[:?Ub7a8QM_g-?FFdd1(e^JR:eY;)FK[FW0\ae&Oe\THHgTc>E<C>R6N.;)JId8
V_CW.EaDd9WA/,PA(/N1S([PDI;#\.d6Z+I_8g1N4#SRU(?L(2KX#4-3ACS/[<E-
J];#c6JQ?Z53+f3]RFLBDQ=/M@(M]KB+)01/#.,+TFg+?#3EJA49T=B,XV=/S=:#
M@=@4K)V9BNP5;DZdUgM1a(-\UV+7FOR93ZdJL=]8ScL2[6G>^/<=++:AcH804@2
9AF8^Rg(?:X415RY]]e07Z4HQ-ZA_P^SJ0Q;4@W8@\2\)^f9+=>-a+>+T^:4E=U?
E6JFb8L8^,J:DIWe;[MAVYag:bR7Wc0R=AZ:LVH5[R:d_8:NI.P21<LO3:EV-(?&
0_F793-eV]E60E&VJ+(&dcRdT2G4;YDR)F[MKAV-;?KF_FCAG.32C4g(_1E1Nb>L
NFQ@S\06ET=QfJ#J.](RE-^f9[5W+V]Y=7^VQWbD@-Ae\7(0J#X5CSD/B\@D;Y.(
]E_KWP<Cce7Pc-bM]FX51:G,HJ05c\cd/APb<TRPBa93[C&MU=T#P3U4D]8>\FH+
L@3c,411Z2Q>4C_OE3d:UeCA\2=@Ma9a8QFdS8XEK^(?3gMA=B,K6/FRAU6)=V9f
\G/CP/<>4NFcS8^TZL_dN.^5Q69]KWe9#.=R1<_79Ra&[S+YgFF\cd#&\g3W&5@\
aARCZHd,_TU^c@5@0VIP0:O,eb@6@5_E[N=J-+=ZV8#AF;H-RGLI?<Z1e/\@T_V2
af9X=LBJ(M,:Sd5_MLdL]_a,DX[C&,L@/71E)U_S:<<0R.c+PFR01g:1-Z=5=CMG
-e:LN/D5WP,M\0J/<BEC0T-@LIQSSKVH;7:DY)b]#M;&\aS68:NU61(TRA:M9(6;
=gYT])a(HN=/836^aL\GL+(AA6Ec,.e>JC@FTA^I.a@G1ABD0ZN29+H/I7K&U2UQ
R1]A#,/Y7+P&GI_5e\TU+T6+);5<QJ>g&:IVY[aXH,H1;L8fNg\+YE/>Q-Y]aE?7
HLMN#.J/BKTZ:?8S9,?W(B>6#F=R3H+,WfLC>dZ/A1I<P9Tf.2>QM_6EKLN5QVF1
F1c:Yc&W2NA,VH77c<2Aa[g9TWV5(<,&7LCR\;&0FE4M;3bQFFMMHVBdOb-b63c=
)D5VaN321UfJ7;gU;I67.2-5fE1?bH+K4UH\cIRL(CaWZJ78dO5N]^KfM^MN[d.E
eV75>ad7&0_\-F[f,)?P@U=333(/MG-,O0H_R(349OEO/E=WaC-PMf+C.4eT+BQ=
e<?4(O\1Kd0ZQQ7S40;84V7]e(:Pca#((\7BCDWaDe_J)=&N35=9W[7KW9@c8+M^
gS\D_)<OKd@_&+1c=FBE.6:[:1I+/.)I#]SGWLUT((CZN.+A6GI+H5JX>c1-^SR.
L7+g/H?+V:AHg901>OGMH7^R&#@+^8H7ZHOOI6(aD90=Lc5>@6(+R;KNIPD2.[ef
58[f8,DK4@:;&#YSEVL7WaaA2MD@WNXIf=>IGJ=FB<\0(EGaDDdV8HQ]#_]HdF@;
aQG>)b#X)WR(c8N5@)\O]CQH]N2_N)T0UL6c4[aAO9_OF:c:cPdDFII^HSB2LEON
WLI9/&M<U7T0MD#P^_T7(8Q]<LFSgdcegS.B@;T2Ab,#V11>9Q?Kc+4D_,?MM/XT
COV&)JN_UM_QgK@FO2-a/C[&=df?f>2ab^QS,LgX4HbKQg-7QXbE#-4GSc>8804I
c.K&eQ:=Z09<Vc<\)MA,80@T,bW#A\0_.=a?M,eXJ-g]9SKL3g;Re:ZP(]KXC0ZQ
M]K=LeT<dGPgeJ4WK+I-D:@<M[DV&RQ5PcQ)/]K=He&J\Z]PTfPFC_PIBg)F/IBF
:KXaKb&AI:=>C]A:[dA+6>W;^-5CZ]O-(fAB+g^//OH\>Hg++Q]#eM+\ZX8b+529
=b684f^-0\T;3T2AH:?54dY13\AMM#;VY>d_N#:[ggR6BC5>>4TK+cG3ON=?TIH,
3Q)>7H\AMgT#?F=VBK=3Xb=ZOMZ@[\aW)O6\,:MF[ZI++68gN+eJcPQgdVUE9I\b
59T.6R/\W@5/c]TR&-&,)a@U-Y&PGSP/M)@RM^SLc0KaVG>\HgGa?a(T#GM)]>dC
.YDVX]D[#N>4@H-RJG[@eVPBW>2^;M6J([TQf?OY1f&W6UN?+L0&&,UTL)gP(_A.
W>,,Ne1HTT_BQ;;dZ2PJ;DgX&42]3\1+N>WDRWS34/J,2V=0[\N]AKEE0VJ=VfgO
-2SK93MA)8TG<f9X?Y\P,?+P23,X.=]V_NQ8T&A0#eIC,+G#f9SbDNYe(&_@cHW:
K/JN2G&.?Y617&>ZWcS;SgC-Y:F+bL2E+</RRRdIMgH+QdG3@O9LIb36MQIe-KPG
3M9[aLCKHWZR1-dXDELa@@=PeZd0cY@U_PfaA8)2B:/J2V)gP/3]/Sg.&EL;?eY5
\M7FER5[/-5REUdM<,YM,DH9Vg4?+WJTfW5@a9P-LJ&MW=ZE2<FeB[(]V_H-SbUQ
D;Q0\G0K-U^TG#>9eSffCR/JZbgYR-VX<<SM8=B#)A1?H>G^DfO;XacbW;g]f&b=
VKBOU)E]U#41?.\3\^XX.Ze(MF#MD+f552/>a.,Q=B[9F^XgYL,geQ(b^F>A]Z>7
I7QY.)VFHM?XU-STb)MT\5bVUFQd-](e-3QP#-4@J<CI=78^-G:d9H->T.71/^O_
\3G.X4@RQb/0ZWJ6&QP>&@>@A]49gJZM.@[^B20U?=ZfD/T<P^g@gDK=N:,3E3Ug
25Pe>7A538&;O0R_\:F^7f-AVP](>8KeTOVW6)F=3#.1O9#?33e)b;0[Nb#ZecY_
].)&+?a3gJcHg>]5GY5SLe65(=N+ELT/21)XY#WK/>5MY4MM:Pg&K<G]/4)A6c3R
Pf.a.VAAU-4@:,\1DE+Q+>&4XcQa,6c;6+37Z/6HORYdJ[:FJWSMdgV294Z0A\Q9
dQO)<)(=-0W\8I)PDZ3c,E^f]-[f(XVH@X:0BDQfY=[:(/9VZ##5/eSDYdWV[Z(6
>B&PZ]N3U)F&gIKVE=T><=8ID5@b9VL4I0_K++^&M+SM:H&\5X@YZ-+I.E\E(=JS
VX,E&WP&b\DS]cSP2OIC[\D^KH-fPR\3-HP2JTMS^Z=5:1:ff@0_8UHMaaQZQXe/
a,2e1cO,]@22b.ReJ9\#R]5/cVEU?/)GZ&R^4K?8+Z7<_SH__CGa/ACI0PQK?0(Y
55C4:_?a50H^,FbZg94f-Y]-GO4FMC]FJ^;4\LR]b:8WLTe8<-aD&cF5ZHVVWcVA
+f<34=9daJDbEA78:#XL+#K);43PB&gL]5P6&?GP-X_59_PJZENgbfRK4SN:@;DB
N95-2I]74ALBK2^_MZ[XB9]fcKa^;-S0U)<)-H[W].=J_Reb/]fIDZ.bWK-K21V<
#HR]^TMXY\WQDfQ+Ve\VKf9D^\Z+a5@)4<Z3a-9.>[4O4f&M0JZ8TH99125HM_VA
dXK0=]RU.J8+D,,QFMF)aR(K7_1XH=-I)/0+KCZ=OMLZ,KH[b#>[STgX[/&SF[e;
,Q1Z-K:#^cHM)PLW7\@S4YSecb\1KWd&VPOMF=,AUMS1Q#:ZEWC_SS8]KBa6[5I,
TbZb3WXY1T3_Da>HJ&>b20P^)T].Q^57NFOM&a+b^M@)eLJ]2bM&;>PZ3X2WU3(+
_a&@Z(YLY?_O@B?&J_4-@c_9.Jd;+5PM5d^^=Y_@bT)H;1JX.TNR1J\ZZAE,DTKX
-gcQgOXNB_IQ&-ga\&V_QS3Kf+#GT[0CY9)R7^]LfC4Q;B6d62fN&_,]5_\5O;.0
4(ONT4WT7#M0I?&S(dUG[841LLPO&\6f8\(^1dN,/&Y)@JH>@@N+bbVDL\IRaN8>
1KK=bO7DM<(<0;P675NCUX5&#^WHDZ1G,cB5+X5FCCg@\W&-..XSY)S5=S6Y6:XM
@]Ua=ga(bI>J188RBY:C=;)YZg&XMB6_@c_;^4O^EPH5[P[XHSd5W>CE\bafFF.[
[##N,KLPeY(GgR)+\Pb\ERXTEg]A)cT1@V>-&2P\_RUI&<,bJC;3)<G0BgCSI5G=
(gE+MRS4HWL>a+4;_C&\<@>I4:I],6YKYaY&2XUR@(4ae+/JN>^4_?@H>8UMKLI0
_]0EXe(<I=EG#cRXTAK;)&CSf5JATa3URNK>B4N\N+0,2,L#+]Pge/KB/D)^bNaR
bSVR0Y?S^1Ld]dG]4L=g.B63PS38K.H_aa:(;2(5&W3Y#BZMI.VH;Qa\C<<W<(Mf
6Z4,._We8M]YPN>(H<bVbY2^7@]@5H[@;FM^>V[45bQ]R^@+bB7dNe6@>MeZBfH4
J709YdG.[eTZT:QEN:MNAcR5:<;HZ/A<fO&^1I?]Sg^X)T;H,W4LeN;bQe\.=AOB
?:JB=PL+^gDa/O_F>2RDZ01OAYV)L7321Y(UKQ[:@2X9:a@QB9eU>YeC_Aa/>(F4
fI<D7_;N2DLYg5<\[NU60J&=7,82<FX#91[/UO@V;>38K2:bB/1PF^^V\?EE;7ed
G+X>>)^^:B??80\4+<Td-O&C8YL0LWaRU\J.@N39)#Z@e@eT^=CBa?ADOaLZN:b-
7WYL)8g[.c:5b,eabU2Z-/_#\07@EF:7ZYfB;?GDd2_H_@.GB7O+TX-Id<0U+eHA
KBC]O,ZPMd)6D@cX-9W2-abO.HgI4JMZa.R7AYUME1KO1CMAGgFOR4FAEP29bgT-
bO\(]dJ2<aY_)1a,@]9I)-3C4/f43EeDbeOP[d;g+.:M?YRb=O1f+1FMJH;I^YAe
JY^7O14fZ:#eSNNSf\E((QLg5-2f;D?f))/B3<B#:(K=QX;/4&\e&KUbWbU;:<Q7
BYc(H0aN_]+/2+5PWHNB0/&D.&9caeJT7N[)f/&2dZ\\(R-IEaFMXd)dUff6(b@#
MNUI.X5d^6S6-RJ0b=M^JG5db:<@?68KV,?@=/C:^aC9?;UZ,a6cdCK<6&:^7X;3
6E]44=_ED5U6.&L9ac4VP=dD<AZcEM=M5B92LV5Sc6ZL0NK:,.>cN@4+?_W^F==2
FFb;bY8\bNDBSV+Z>f&+PPUdUT4;/8CDaWMLTY]LFSeB_092EFPP.E_aP#^97XLN
X-45S.dB&9[\QSb+2Y@BUK=?UHRX_d60\)7fYFO0VRa15GH\LI)]RS0fXCFY?W^)
\GfF#Q3.;GLIAR1#Y0P4P00BRI@@E6@M3[RG3Uf#Mbb#9G)^X=:@))@BA_2[M4_@
7##\IfF\bKWWK_L+&R3VX?g/D2=8&:cS.]AA[QNV2/Xe,3ASHCH#I\CbYLUB/QZ]
YVG<b9=PK1,AHM4/R-;T5<03IOUIAZ=Y[(-(D5BV)>MCWeVRb6NGC?<M[J5GYG5H
RCHF)Z3#W^S-PYO.4bB4]FRKD3L<5R,Q3959.\Z-,DS(Ob^aP7e_X,,FM>#YG#Db
99b[&5-F&e>#bFN]aHZ9H6<W8C?R))AeML/J6XFC7;C]S1;K.QIa7Qa:D/L\ea4^
&]WZZNKdeP^NU7U9H/Q[M4&.Q)cU3I2P26b0c3RRZ;-ICQDFZOQNQ@f^)P)P^,]Z
=GLF;=&7aW[\<d)e?^@/S@?4>4C47LcG7#Ifcbg.f5VL8;We+KFaN9)MPV(bPga7
0IGTc7[,3_V4U7:LN1\SAb;C-?1)^>B:Od[G7B1gK:4C,3>C(RYI_+fB?X:3\VJ^
X+?X\XILI6:b@b_.PT79\P^/H^^P?1ab#\(46(T^JOcL?M=)DD@_&0gY&GE;9/Q>
?UUR.;g1UW87)@#f72:NS>B[L?cI^_MNZ@Y7B4N.NKR39HTf4=,9JJF_QT<Pe+AB
IcTIL@7)?/_PFL(<bUT63N966DJ@V1WGS.+<f>H-BC+N;TdSB_,aW(4(?B1eeaU5
7]>@gXWG:_)Yg>Z,QOW4,R3V.fEMOV(b1P^cM1O>HE+-KR)AIPK#Mf(,Nda=4L>U
7cO:GbNA?^W4L[X5L48_M;^-fIGJW^GR7^(RSR673FS[.I^UL8;=/42L+DPPW?B;
HW#LYDa:_Q^2AJMP-2LTgGYQZJ+V1W1LTB:;/(:,LJD((>+g@0>V_BD4>c)cd&:I
8cSBRQ&g1;QZM\ZE_9KFB6W(0)g6/-N=c[KIe])a,;3^M@YZH4#;_eGB/AL60B([
K&Z^2Xf2:O(LO^c&SDLMMfAd26DX=E0+=06_;0RFf]0WQO/LN_KYC<g,(ae4,Z91
P9.6KL/#U9a\e7@.NN^SGY^,<fSJ?e?4X_0D6B(VJ/1E]HI]LCQQX:?418<JGJI_
R-g?eEVLfeWQC/>-Q64BQCg_//@2F830:[_66:_c-[X<X6\]FX\4>+0_LV7,]^bG
L.<,18SJAZ<9,SN;55,L,>,4Z-]CR3\A/8W]Fa:)@Y-Ad#[;=F#IM35=?b1QWI69
M]X64bOSSE^0O1:,\U0^5)B\\f-BME2)U6ASDJQVeZH#-1)SQ)2S4<E30]+BOKc]
[UP#ZX_4Q?#ED99R3\:T3^K@>/THRMUCVNeN#I8M_-ANd/W5X3a\O#XW[>XefDd[
daD,0:H@/[)4f1IPRN>&d[T<55_Q;A/aHPZ;ZPaFJ/MH/AbQE)&IQ1g?)1W@c<gM
XSQYe_?]Tc-TG1XV8>fJ3(+I8ZVUeC1IR2UbIS3P4f75GN;,.>D5daUKF>4>ab#a
M\0Y9];1S&WM4HWKY&E[R3AD)&ddQbP?C9a.61<&X?2U3ON\L(:1TQ6&)/:4fA:Q
.I)<<X\[YF?4c3\2V(8)LcV;MADLA4QGZ&;MNH=)<W0O1FYDEa:->+aMZZG[gILa
e3SXM#N/ea6fS\Y,M,QAaD6;;WAEb#V8#I&T,bf</.PBa,f50)R?^Y_ZXd=L7O<Z
H\KL0(H+U)+=9@N?YD7-Y=VcG)gX@>FeJgg5V1Yb87.;5GHY()a1G[@DQDRQ9>S9
X7eW:GC1>gbP7KQ]T--5bQSJ[WFWJY89?QH@HC8T]N@;JZ)GgG/?I93&M[Af?E&;
W3]4C3-]N=@e:+S<)(^2P?CY9;YAeCSR/2D9:(-6DK,fV+\D]KB@#@@JA-T4R+\,
+YR2RX#Ff:cK#PS=A<9T.d+_;09d@FOBE&.>&\C(6>>3.O)H^d>.#VcET>10#KA<
T-V46XJXS+FSg3Sb,.^\J-_O-E59MX[A8CW.C2EJ;BK?Z8K1CIKQ1->]075GTHG1
ZVa3AGg26_?A6K[BNO:3Ab>-]QTD4R8a(>+beZf7_#d8Ed<);AH0b52>4@/gBD@:
HI&2(J2bHRV/TOLO9RPb?Cd>0&L2<J3?Q+PZ:;H1]9De]/5+PWY&3NH&.X7H1QL.
:\S(VPA,F41SZHVD4^@dT:?W1<aR4a(^VUOS,:G+LI,+H8IHHa]agLV\9QJaWC->
H>DDA]8?52KVW.1/.)ec-;gD^AJKO3VGMRW=OfFb1P6(R.U+:3df[Y/KP;]JRCV9
_D&?\L1TJA58g^(RMJ>)Ub(9RT/(gJ;aX]SA0Nd-^#^[O:K^a)I.ZSUFU]R2b;Q\
<QRDTK0[65V;Ie\2c?A[K0L-\M>KK^A6_I5dQg(.abS]ddQM>FLVJO)>Ce._3da8
\^EI^8=2)F&,T3,\,<M?9[\3<+]UEB(:?64UTAVLZN^e^d->8PPb\2PHa1V?XOAd
,gC:2M3D6/.RQ&d7)4.?7],VKg6<BfXURReFS8Ke7],^)&E?4M2F2cF4Se4MI/4K
Q-5e;cA50-,HbPU(&d89?:XbH<WV8fS0DI<U9&=<\bEIaS4HB-OOeNO(@Qb39Q<G
)I?0:N+84@6BFK@I65Z(DB>[;19+PFDbYKb/2XONd/NS[[B)WE(;OVRaXD:>KE&&
EUOaG+bXEgQB#H/ZGY1,ZZ;_EJ0HYY44?#L=71AR)fFY0KSSaA,3_&aC9D-.B7.d
0f/^56T-XVS0Bfc2HKJOJHF7/;AU7d1UK[X^P#QY,[DPe/BGfI&6/B7Z84SIZS6a
ePBA<316LHX6O#-693G@;.dQWPB7N?5Y,YB8VQXM-&^.]0IC40,CK0+[-<f/4S4:
5Z]>Cd3I-=[eKHR[.F<9T/L^Mf=Oe6b.M8@TG>Q:=fU]>8N0VR6BY6/[W(WPeNL6
5(BZ+R)F3aIe&Wg2T/?>9Scdb&2c4R)7O;T1;A-\9W;B3ZYP4:1)R[b13U?P(Y)6
[B.YeBXgdHG_.ae<K;eA>:UD(-Z^.9OLE>K/<EC9D\P.[)]CQC(\ObVS8UJNID8G
B1VW2=&3#>E2@D0N-[?PXcIW]-g41\8FFAP26d;^8U)N/]fWBS3cgRB</5#Sf+0#
9?20S>]0F^=D5PPF7EFTYHT(@1ZSdcdS)d/eN=4\6YU:7+5Z#,J6##9J;S8=/#EO
bI2Xc_6e:[SKZNV]/C;\T>K_a1TQRIWc/Ef[J(,O:Raa15^[\R,5M1XVY4)5NRB&
JVLI)VW:,f:CL?EH?eO3]1_R?XcH-_3?)^M[UD=)+LD)Nc)N?FZ)F(cYZ-3.c>f/
c)5?\Nf@XaDF_Y/Ja<A+#DIWYgKB5;E/@@e3[,YXA;gPP\C&_bZ+.N_)7,f]?A<I
H._BZKD+1D.W3HTJQ3G#aM>a[KaWbTU9F6Fa;9D5Z/#[>;<UbQ3II^](0dL2OFd8
3VH9@C.EZ]Q@Qf#6f@O>b9FaRSM-7#+,0@;L/I/&CJ]<d7G#W^#2c;g@7RN&B@ZT
Pe\H11;&?N-B2CJS9.a4_f<\,?<D72[@.,b/PGDd#>#1O.6\dPJHI1Qc.fIgA9U[
P:R&5]39L,3DY19)+>/D)b#I5e(XbJ-57)CYFGPL&0&W5/=R0FQ59H1=:1U#b_B7
/+^BD)4e?ZWRVG]]9E1=);H(b9;<#-Z)\6S[c/N0F7O_<M]H\=)XZPQeCPG_1<e/
5_IW2[(2K/18LT^Ne5;PP@cXV]Q],-aDc[0;T;\e++>D4#KPb=.R21V-.R:0-Y7K
f.42+=Ed:JM)X3E\K+69S<31I:DeK7JLAG:RKB]CMZI>4_9eN)d=IQdT28;7g6AL
JHb;Y3IfC2^NV[N&bQIUZ+R<A0C)<8?,F@ZK<YHK53bOC1C3&Ra_OQR7Q]&J]dEV
&HV=/UaF6A;HIGN@84Y]CTS>,3Q[ZZ?UZ1PA6aMWDR#XV<_#H#:61;0N<IUHM\WA
E,70VK-91M;Sf(TZ#^3cYN2OaLAaV9^>,2JKd(-H.EE;.7#1@G<4H(>?/X<+)2-(
82<KJ2Nb+Q?-F@2U,#dASQFQ:K.Y/Q/NL0SU&[IcCX@Y+8a1D^>&W[].))WDH04;
d(NgVD?#\cCgZ1;U\SZ+V@IIHOPK[.6Vg2OU23Z2;)XgJPUe?/Jd7_Eg]UZ,J5D6
B<g\8YP80f>F:4H6R&e)-EMYVL(\0b-HI510,^_C+<@\fffN_VI)g&/IT:Gad6B7
E),3(6:QbE,9[]12YX.]]D,g@PN&^?;,Ng=4SEOO7?3fT-7\?Vfg11>)+\,XRDO<
e3CS6g,MbfQINZ_5\W&#3MaMb943+;BNY@UK9Q]dS\VI+QI]:9,UfG\a=+3:S+X3
_ZV2VWT@VAP56Z28BY-3[DFgPgDHOR5#G7\5WO1FcOKSR5MYP/<BH]U(VFN+Y264
_#U)_)OTfgQ-d7\QPBV_C&L5&FU3IUf0V5F)<8>FKZ]0-:#g_M>85X\NQQ_g-1.,
JN2JF93V^f;&I1E\];[FC+>C5645<_1?9HOW+]4DYZc81&IUaM6>>G/+BgHC+CNY
cF,PN)PKZ(d8FZ]T_F[@(E#.;?(I##T2^Zd02S1B_:7cY(GARK;IKOVa.-4EZ4Rf
NEZJ]OA@3YB=L7Rd1]N_<CeXG<SJV<0US)#=VTa_a85UPYQ3\d-Q1B8PY&33QO5-
aV[][>>KCH5]faHgXbED4-OMR,VS]-6\O.://9X9F0VTQ#+0N3VIb^G\cYU0(?EM
<2:aE(=:QI8)[_\TI0@0c)<N6>9I/ccF)B&V_^\UAVCMOQ?W7WL3F3ecCK+2@>a2
/NDT:Lf(23P#?YB>@g#H-26IRN>1T=+:c:BONF7C8)c>&c^#2U)L@&-8D)R>CY1L
:C)ed#;1XMEVB82THA:Q@+-ZIYR8M@WcW6DBDCK;]18SP_Tg]/<59gR3AaeD2cHW
Q:4eY099G+PD<<VI5+NH6WY:fISHLQ0+Hc,]<@MIM(6U+KMLA\T5/WVWH\Z@X(A/
\RJ>?Y^<@O2NGI+=&f/;3KF,;3^AHPUf[@e73dJ-bbFY0:-=01BJ,\3J@e2<6J)J
gfB<EP33PSO\QL_VbVDdd,0dg;)DP1WF(QX3</J/MLHMQG1HI[cWB96V4-^(](gD
[^MS=)529.?ed05Fg8&&6\FU<:0fdP]J>dI,92@&fDA4QMS+S;U#8Z>,MLGM/8]O
6-EXIB(<Zg4(EKL?c&9+A0_<3YN:YIB=R.>-M_GU:MFd/HMO6@e.-/>W&f)T[:DP
^dDdgO+D+,RQZ/ZWHWD=]-@H9&:_?&dX,H_(\JUZ1(@V;gTD;[T5Ob.daR8QRN?N
DZfbNG&0IHM35_N.J5@\FR&_gZcQS]19\OA7.]OW&cN^K\[eA01],NHKF(bB7-g5
4JIHVP([AX5Pae<R4N:/5?#M]@3>d6C.QdOd[+XKP(3<Vc],N1#1_@:1.WNWa&6+
YBE.TKCDXW:2;IJ1CEX#g7\T0T9RL4gX\:A2,W>/Q++&&0b)gGLNRIK:K2e.f#+8
6=8C;4EgGM3[WUg+>-#d_Z4@KF\/8agb1<>M<#WT[72_IZ8(^1e-ad[YHUfZeK?e
=29/a.<.]PC._7K55T_Y0c/Y=7?^FU2=:[ES_a:]/-@UJ47[2a]SG5\<a&^F:g@8
<Z[HHWA0GCD:-DN7Ba=KFB[5R+.<>^E06HPaC@X/F;NMSE;?-LaWTGE:g2LO^V4)
#VPE8S451&2eW&a?)aW;Y1++<>+fV4[a/@(9+Zeg/RK9[C.>19aV4@fUD1Ea/0GF
(#CBT+99+(GeM?ePRT^M)b[cJSRP>G^@Z7@VX^\f/H(02cc[OU3baQN38]JVH:=/
X,SbgKCVYMb513O&82AE>eD-W6#Q#&+0K_EYBc4&D/1G^+M_N?2@>>&@:59Y\J/@
LG3P-c,73;cPRb+ALcE8#eY;[OgYZOI(_4EFdS3e.Y];:T+9GEGR_8C0RGI^0WBZ
11^ab[aJ<-&(H[M-SMe4e3.4:Q\191c8b.a_B?KA2U6XP-(0=1#63G[^2;0><[>+
2dg/NEWW)W;-42+/I?5^2H,862UgZe3DaccXTM5I@CMWA5C@,CRM;2XH5WbH?>RT
,5C7.=Rg#fd0fOXedb0N2C_8/XCC=>YbWL+K@M=1M\HS\N/<IQK<QC6_M-[V,G#F
Tf55d&==N(M+SMVS^9#6?+SL.T#0:)#>+2K2O[dJ]BeASE)&Ga^SXEHQ-4=6c2O9
]8<O3gb(8P,X)?ARS<M:-DaSg#\W2/F51:4G[N/AXUQ,^;TdaA-KM,b=M?F[#-+a
8aLCF8RAg?E\RI&.+8)5?^/)96:HcZg9F+Q7VMc_-D)6K1d=HJ&HZ9e]QV.>18W=
aQcd/X(\OMO#V/6XO#:P@]eF(P3H#8:KJOgU4V9DT/0L6@BAd5\LPe^06T)BK\SI
EIGP0d(BEbG#[M7]GVD(;JA05OBb\b@b94_FJLWU1AZ8[B&.]D:8P(.TNaEbUIM>
^g0]90>#&SY07QdF,SCZBL-3fgC97CZ9d5<<.M]JL8BJ4f(\gaG.Qb\-^G61W8E\
2Xa[(UEf-_EW+\LSFWX1(/+TbFN,.J@4CHK5N^F1)))E)-^-,:16QfEg7?I9JL4O
^&G3<DJ,7P41V<BZ6(d,U5>\GL:F(NP,AaM=M@R,0T/#M_.YO\DMYg\#0YG3URS5
Q6dg1E+HRUG#caXC5LJVSbOV4^cR(K58C7,79f<K>[I?8-NbY6(I1QL@(La3FV5g
5BF[[?2MY\GH:&\eC1WfA\M<@W<]2e+N\K&5C_D6_I&-P5?8-DUa0Ve^P2AXW:(A
CEBD&3,C3X4HA=_95_BHD@/OKGGLa8Y3b=BWe/ZB/6TVf:2-gcP.9[-Wf^\VY#5)
[NP@b<f@5dUA.b#N2Q(2HNKEA5^0]2X-Q#QKC?b@XaBR.QW)Pf?7(M_6R8EA1@Wd
R-V&67Z;<c9B9=9R6)IWD27LAFE[4b4SF9eUW7#I=&WW;?bf<aXf<@_H<b;g-8cH
+F?HPeS)fX)\EI/&+<4I;K9G9O.b\>OLETf7=WAL+J,Y+2/+<dC9@fN_F7^3.V)e
O_]M9EI=2(65OXPJ35B]&AR045K2HJe<1FL[-gF:HZ?A#]2+ENK_,URVSf:W-6:L
U\^2P+RY]+D2\IJGe1J53@>f@f](I=2CM7P#7_E0R2Ufg;OFd1&#\8ZFDd_@3QPG
QRRc1[:;:DdU9#O99beYSSK.50#WVGfSXTULQ-&[Sf)JGE)1S/8Z@@[@gC0LR??@
D&2d@D@QgN(BF9DGILF(16X>&c=aA+.fEe#9ed+-dH/_R/bM)US6P[bMfFJ+)>;;
91E_a=EBCK<?)DK-+[J85>-Id-Id+]9J,;9LWJO^8QQDgafVV:De[G;T,)^J)[7>
LU_AGD>f2:XA9V.@bAG;:\.Sb96Y)IdDP#+,TL9F6=Ab21eCGeLRX?W_bIR;H@_]
\MA?.WIfSTKCTFgfS+fAU(5]K@0MH8H+QL8fcTC04#6+Bb7P8U2/GY>8_^ANMCI;
IEE#MUIba+IW<FQ?FDD.dBE&3c3+\7M5HB(A@D.dFT3/@FMBRf_:(F&+B@3+RaC/
_YY)50L+)V_gag:;D7<BaE<L5#(fY&Q[9V@OgNX;#IH/35H80ABgcLS3N/&#U[Z2
Ia_:\3gB:50IPRG6B;CP)Mb\906N/9BA>FM(2#6S5B:cPET]fC0=_C[e,=&?B97A
TPa8&T-&W:bPL0W;P1]^(I.@W0DO,VZRH#)S&71Q(7;#Ada#1)K<D(<[YS@G?I]J
F_8Yc#ed>;7(P.6U@SC8Gf[@e01,=E7?5\WUL4;b+dFYR^V&QO]0eSJJNd_A?])H
7b&6[9aYDY+/4_E)a4X[:0d+1/=.Z<_3aY[F7+.:>AY394@X4?]Z0MJ)>+0/YL0d
_:8I36@J+cDMcfTY)6S(TAZ-b-GJ>FC?=W3G,DeJ@=g]1ZaI^#H38feaa^W-4(Q+
2I]?9:E#W^OQc):)f4J0YEA_]-B-De\1#(9,@CIaa=3XJ<B;K[MVWI>gO380dE5P
+e)cXNL:8=2Q(D)^?7O<:Q2U82G^EZ>-7PIJI.:GXd6A@Y3+Q[9@-JJg#O&Vbf@N
O0/=aW<D8a<ME;K<O5cF_2P1[OSW154PTI[;QM#R<]#O\QDQ-,FC7Q,(J/;OJV0)
:[UG.)PL#(5O<I53eDD+ef?UFDRHFXg3:@DO[KK3G9<&Z#KFZ]be^a-MU<4O1^R\
Z.Jg]Z<g+Gd]^\=AdAX=6FRSCb0SZ<cPKFRA:/]?;(?LJ]BZHCI<ML.8;]a-<=HY
&EU6.^XAbQGJ4;]2gM)UR^S=4+aMTa-(7+dG<]K#Q@#:/e1U?cJMRb1:NC0:e3NV
b\#H]]T#646\CM2P_.U6@a5S6T#b=R]2LV+,>\g#IP;_/0MUS_R0&7R)9@\gM[<4
<J&+WD\b8+P77F077S4CH8B#V>VP-Df?a5B?\+7&_,1>bH>G[X93>GfE(\#//WH5
\Qb0P4:M)egU1?FXP5J13^>aQ1LE2FXM-\=Q]QC=/9@MeH;ddG@O#W]NNA(=_2gB
21eSL.AEdA5H_;4JcRHYMU,K5W]E=Z6YgY1OPJ)@Ad\CN#d5@98E;+23-QNUXY\,
^2,9IbJPcg+-:VJX.aS0];-R[?WUF^346a)7a??E#&7GEW5T]ID\J\:c9geO\2^4
DBT-06^-6EeHPSKa56b<eHQdAI1L#?V[-]]e]@07MdWGM38\>dG)6=8W+I;)@<^a
1N+HXMK(8D\]\)[><V2QJAMELNV=\dH>FC99#AU,J-SG.b^L6_d_T/fDSSd]/Ddb
3K<NYZf[F:Z?5VRKT]^JEWMK22C-Ng=7H@C8^LZ[L]];?&=+YBUYI;(0Wa06N5\H
c,/Ng\#_2V)0.-6YG^A8-dAR)Pg9V35a<4+#JP=8XafZA1VUb\+0\\KKI;F3EIQ3
N^fBCcM-PJ,?d[9T2@7LE5,PeRM_CG@eS[#O,JAR9G2CGCH?\M-Qd?bL:X/YY+)B
W_7\[5Y:UT+L7J&X.Q?c0+5EQaQ=11I_a?0cQH.dK7&7@GbTa^CRRe#VA6O=;M&V
,Nf-Z).8,;.0.YX,PbRLQc188R]ENL-\<)(<Pba+&U]f1?A<CbILT,/>CEAJ(.Ff
g=<e-7d&^FE-_<^)g_bG-,J4=WT5F73^R+I5d,B:(A8[==16UTgP\)I@/_DL5NX2
_(,XJ;cL5@VPJS4@27F95.@RYJT]:cO6J=#[YV4U[DK(K:4#f@G=OP@OQ:M>DQ3B
4O<&@8PYV40^8B=E,BO:P[)J,S1F..9PI3VCCgKKe1Lgcc1?b]<._8^BA.1[2b(F
/3X1;[Efb2[=_MU[8+(IR0A;[#RPBdZ2?&fLO7AXIGba^/\Z9((Ue;(@a><DCDNJ
GYI1UCV>3@KA#V^X,?P2EB6G;[.2?@_4FZEYMCM\288g)6&3,4dAg7V.LDg(>Y?7
WU<_9R[<G=S->VO3KZbRD\^7?d1PVBY;HSYH=?A\+W3F>,>?YG+W^57T?I.0c6?T
-W&1O[C^S,H8eb)OM@4UK0P.^UHbH4;7UP=&@U:<6J;gLOH?PKU/2>(C;Q.PDH[2
Y7QMZ,F\)a-WFNI\I&E1(g9&Tc51VFA50/P?_bF\1)@V^)#F,c.D-a;_:&B7:/_5
#ACX.[Da]aFH15;,4c,FCS=7-]bgA[-LY3DM56[F)^-6?V(=3DRIB;W:I1/:W(N5
875[YRbY]-1?E2#[(3be.1Jdg/O9Ae.Y<_?\=MCe@W2.eaE-U>e]DZ#B(Xa#D4K<
g43P^GN3C:Gc2><T/1]G[R9BI^)./SXBbXa(^QTAG+8]IJf&2aJM+Y4g89I1Nd1=
TW1,=\HD/fF?TVY1_b,8V_?AVTB&Nd-RJR0NY?7P33L-BINP=RVM-@_)RJ,S<.f/
,(RX3)[a1H9=DV:+;F]^+)cQ#NZ;@O8dZ#5dZV]8Wf.0+K1WdU.T:?6aGQU>>dW/
a-cFN02BD(R@(eA@bTNMA(aW5Cb>C1KJ>(OO88P6b1A3PWP>NDT1<U][O5g(UgCQ
+KHT7\[GQI6-7TN-8[bR56,)=9J(7a7O65c66:bMN9Uf)/^-D^V=@@&c=I[@c?^8
#[I_3^=#U#IP8,Y^CR\UTA.63S;fIf8DO#MNUF#-5d)_,F9#&Q@ZVcT#AOYODZQ1
:aK&f?ON;I=a>[7eV/\Iba6F?fRP2I0=eZV0CW2YeCf?MU++MfPUgggV7Mdf=93+
[&][[Gfc_KHgT5?eU,JZ(EbFC7L3)^/7@GgaC>N@VbAX-5_&-b@:@I/O<CE#4]ZI
EQQT\GN.Q_)McOMXS_WN1/B4D29Z7L39Z+d5LeB3OZBecUKgHRYB-L&86DIbDf<.
);2B]X&f6X4d:c==2\\RRE,OeH27bI7M9G7PS+dV^Ia1_;@I7),,D0ANe(g6Y/]@
eJbD;+a^+AV?\/<2?M3_?/?K<&;Y:XEG60>@/UC9M0#C:W.?6]I_@2D\eV\dDY1,
P^KSL-,C/HK+&,1>C?]2cF?BE&C@NCdRgg3+:M;^R9=61.#H+;@)V[9bPdVeEK7L
TDT/=a:R&D(>b(630XZ;\<TJYc.WV#0[aEHGHIP[8CS:=]OgbB.b[A(T/K<+<63L
=+0=gUAHR4e&S(^7IYLdU4e@aG\ROg#?L.O0?WZ8:df)^SINGO=7_4[LQFEZT)+T
]1;GMaB4ga-7E#C(G2:<+HN-RG\;7SLK6FQ_ACG2[A_e)f5D,9JW:^+31.;SJ9f<
(WO)-IX.K/NXPB=<,R#HF5Z]gWS<T-.OV?&0=>-gF6MUF2>U.@NR_1Ib.=B7ae>&
8HeI2-W@+&N3WI?>-bW;>9X/aEeb:\agKHV94O[,b?D@TAgBaZ[aEOMV<+@F\0)T
XUW0;/PTD03J2-9<9ACg.CdQIAKc@CO)ID:-3dS_FTC_VXe<SE)MJN7KK7&MX8Af
@,]\#X(C_3NGVX->QPS7C4C4T&<R4FI5@Lcg=[?/+c0VO<:_NRWMW_+M[76(]5)_
R^1)[7_>>81.+[GfS&gMe6D#ZW#DR:8,Bfe/I,a<EF8b1A23S7fN2H+Z2L=6Z^B#
D8c>PQF9P(J)AWO;B#MB:XSG.L>R4^Q3PfDgB.?=bgM0RT0?-PeXMb\OURQ#<:,I
5CDFRO)+bUYQ8@\&?)1NQ;bBPJ01L[UJGOLCDFR3C3<JKXLYU2+Y46-X]7&C4&Ag
R.:gRXaEHe=fJ[7NN5/6^afW\?N)B?8@@F07P5^a1O:)#/3VP^Q,g>S4JU>L7_ba
8NOS5LbM?H9;g-J2DA=7f2W<#[e7ab^#^[]SOW+/;A-:ZBG<N;+0ESICPC6XETc.
gUC-1\DEaW0IP0_;(JR/79c2PA8GbI&3-7Kag26e@O^7g.^,SHW//X^Z3c4HGF[0
LJNR+6_DOOI42HO1[bGc9-)3dDa@0X5[KQ>a;WP<L=0(RVc6C@Q>)H.dYOf&A=HX
M/J>ZG5O3IWIAL^LAP:J/T(>>]V_MGC\UU6GR7:(?B@4BWd4#@I(Z<(9K8dR5G.7
=.0KMZW]C+X>A>c\&H^2R:b=LRZ@cW\^-QKKTec77J(<Qe-CXR^\B)U62GH(\1R<
H-P-MU#KV[\\d@d0a9HKP1c?)OY:+@A<P@VEKVSP,bB[E>+2\:(4,f=f,)bPW#BG
10RFbTI5\g3CL&OO7TO@OKK+_>@=G^D)F7UTZV4\Y2#Cc_,4&&)6/8dL.daH3c^\
YaVZGF\Q5NWYMfNW;KG1FS29[]C(b4R>NROVeBED)R.g]2T8/[GgNB#Vg=3UJ_5G
=[)=/e,8:/AH9V2@G_,OQ2eH)_85MP,1&R).683<5db.FG997>L56FH:b1>dUdMQ
O.1N4f[J07_e=#:Uc:(+0(/0[K>Lf0K:_DE,(6PHcc#DJGc?;HcQ\C1#5IT_eN.@
_<cV7FE0c_]4&#QFTIW<+75_a.9P(Y38bSD9-S_BX<YTf@/:09_SS=V9N6UX@.5H
I7,E@\Cg0E]:(Y9f]@[Nb\V0N-DfQML4THMIJNF2fWe^:7#d7[DK70]6P5=O^VaG
Zb011U6JJFCeeJbNOEN>[AbQKXRV>38b8XE3\P]8,ePM4BD4dgO2a@FER^[-9Y.4
J5^(g4ZCY?AE9^JOMWe,ODf)NA=VbA]RZP.Me9MYW?-;#A@^G@]I?H^J225@d+#)
5S]QFV0?P:CX[J?;S_54&bL6>f]?RRUOOF3.<@GaH2==<#AHB+K3(=[;VUOC5CU<
?E\[cA9NB<;U>((AB=]+A?>9THDDB,I.T9HCBE<V/fCTDgIKd,K7K_B7_7#=[d4,
F\5-_U<O@T]bCBHE3c#.6-_.N>:EVg.^=P5.&MSd&L#7c(\CN,R97Xdf2e0?H:VX
#P,X):cE>fAE6Ca_891H,8PeX@aZ-Cb183A3P9YNKP]7XHVE0Q2WKbbN)BGV0P;>
PI/F=dIH46S8HI:H:F]01&&<eTO=TQcVb?>?\5TfZ7Y5N:I&+&LO1\YF:-;IL/<^
\>R,.[PBBG?1EM^,C0?JF#<CD]V&c8B+EVDdH[[F>XLH98D2@Z^/5YNeK9@F>P6.
I;(HQKM5PKGV]<FfH.K,PXJZ^?WJ3V\YC\&B,>MP7aeW/d;TZ:9K^5OOZd+DZ;F(
dgH?C&ebc;b4YK#2)5=P8f>PN_4N4/XBI0H<YcEH4L)CFTVX@faP3e+<[B3UU+QE
dIT0+f3d?G40:,/FL_f7&]8b+:bMf,HIFPd<\UAO1d->&Q;-0LFaW9>Qf4#0a<[_
M_+H?U/-_PP2>[_F18D3.,OL<XL>J70MH/B/2CM566^#+>^bORB9_eJZR6D/(240
9W&ZS]_aS>bP.KI/H#)#6]T,gb/1M25gJD#G=])A,&JB1I_1H9[[FMH[e,M6QG\-
7]S-H?\HS,9@ZZCg&Q=#@7/.2f96(.WM;ZdNFD=&]/Y#2TSdEZD+?BD21;D8&2=6
F;BGVEC4LLYZ?2,(X&W6:)cR?>Z]PKdDe&PH#[]TQ3b#ed:X@W.cYcB&<6C+a,@c
KKQ(8WU5Te[;J/c8T:0OgH-UV&Qa>FX=ZU33bF&USPIMH-ZgK3@6JOacJXBD/:)9
Kg6F3-XLMLQQ&EG,J]6>710^T/Y?+XYQF([QQ8((JLT?8ET^/=N[V)SDgV;X25FV
Z/0BZ64#<[J4QSaM]><CcG()7X[^]_W;\\BZ7<U8H_2[DNR[P\A=3\TfEF#5dg\H
S9I^a--3PeCS]S3D@XDfB3Z=GXOVDWQ^@JR/cg>>Ce[2cf7H(1L@gVf.;2:fS@>?
]RIHV3PN-:>:J0;^bdGgd(Tc_7H,@?DC#ID_(J_g@=Q5EI,7c=0Q/62OENLYf][]
IMB[VX[P/1C>a9Sfb&_3(f)]WG3>#:?I3]3L7bZAI1AI44GV:eOH6Ta4caHI7)aT
?(AfcfdTG=3,7I27E;YPaD>b+\S:<3<2Bb-5a9T[/IZWc1M7/Z1(]EAD[FbNT?-?
8D0G4Q?CGVfG@U/7^WJ2Ia[Z,>VMEOJ<#)4Q6<Q_YIRC6D=,^O3V0Xe23VYXdZZf
:ZfZ0c1f0&UUBD4Ba#BG2TPLU\GG(&867ZD>O\962PH8P;K:1,M8:e2O6Ib_/c:P
&X7UN]dYW0#G>c&Q3b-@HMGNHKS]5a_:#H;LZHY3(M=f+eNK0A;e[dE^.&;Zb@RW
[??Z\UD28ea:&UN6QR&[O7aUI^-a^C=2NZ0MH#f0I^>9KGV.f_XbJT0/4X3AggZJ
,NH.3D#b@O71U.,DUe3G-=^LQYPGQ+&&eOKF787^B<RLYD&6Jc?B9-X4.X.(SA4)
)@[YgRag<>NA.TVU<)aGIN8fMf:-AW;VU;4[,CAF:IODTF/EK@AYS8RLHF79?aEQ
&E.5#0R+:CZMe?HVRG.gUcS93,]bK1]8_LK;VAVGPI9E<O6R<d(d6K,.4O1]3IbK
&bK<[X55SC>+CGPF<d[0\H47FPUB70b@(GNE:;?Gc2TL\3\g\e0;7QfJ+BOAN\DG
9\O=@;-T?>E(W?JBBONE,,3,]gb9GX5bgdDgaV/X_:FcQb(><4RWBAYF@OdI0@_8
&Z6DB#QK<+^040S<(TP[6^=cISC>-=LDab(S[M@ITVVX&:df,d)Gf:9EXgX2;Z\@
:DB&\-0cOUF58Ye>cH^eM_5<]_S4-[e8?[J6?GYQH2G_HZC#,aI:CL,2#ADTZP;M
2@:d:\\[WPf,1e6.<:9K.,C<-U0D#SLBJUESCO3LY=HSP)\b5gMW=(01J&B#ObRK
P<c[E(<.HUBRg.ZgHdHRKTbO\:Tf8VXTLc&NO3#eTeAPQ8J(87:+Y+\L@FgI@NHS
H+7MC=HN,WLY/(.@8+5>eF5^&=0=C50SC=YFAWP+961G;P:,-C[>^T]Lf72SFK&#
9E@^01:d_g^]A:)LYE=Ea@]-aYO[TFG:Ua7dd[XZfa\PJb)c7>8DD3R92<+O3>3?
W(U7ceBUEFYAJS:1NHF9(ELW[0&:NfP&PTbMJ)IeDJg52VWAVS?Z]^,,9NWZ0MAO
gg7^FH-X#d4L#KD9VabfF?,5X<37W.X871E079\6;H(4Zf31>@9)9OA0^Qd?B?Y^
LFAf3=T<S0WbMHTQ)7U//NI0J0O(VDJ_=BA1fF]V7B_JAc7/WBI;:],6<CGFUVB]
HYD93[SN<2?-251_[<KD:Y;(aNMf)-9.9Hb)cRGb+#GeaCBW:J[D2LP]71.KL]g=
)6ZL-.L6N/,EWCK(ZXXb)EGZFe.2SK0f.IC2>(Zd[3;e<<Q9,+CGR@<cSPQG=O-)
UXO[.][<bd[S#O4];#@b8c42-\)b=FP)TS68S?-]U^,<#f&Qe^BU/FZT^QO/B:f?
/[8OQQ^1,H0(:BV]/cLb#RWJBc2H=N9_TTSg.0,IXR7.8CLgC70>^](0e5P=GIfR
3a>d8R]0U8@A+4_VN;@2VI1bWFAZL+,.D6.;#F82,&8D;882gA^FbQS6JP7+JdDT
B)ab4:A-0,OIUgeFdG1WQ;FQdgb<&/NIM0--)acedEF0?EN[J22C-9HS:28@0,>T
M;8&GTXG,69#NGdgJaDdKTa/c^=]eU0OP00/U)bV\G+&#[Gaf][9F>2-Y[7bKS#g
1&/7682g#QT<)3_E0BF1]6Pa9E;>?V)0R74S_8S[eS;T@ed(@)?<Ic(+71c,I,_J
GZeaNZ_\TSZcT8@,c?cQA:B9MJb3SB?GJNHM7J2K=O(/G79[gWOa:&+:,[;aJF@R
_MHYZ(FB\B9A:)^VWeLM\8bRMeFCJ)b@7BR8R_S&4<-gV&0VQJKa4E(=:f3/Y(M=
?[W)ecT[Tb0[C#,Sc\KIWeS5Hf2Q6ZP3KUFIG]56?K4@D+U[5Ne)(X_]]VG.5Hc?
:,+:SF.WEB7->,L/_//6/-&0E@U]99N0@?&LZ2gM:.L1HQ+@6LML;eH^9XY\212P
+OBH)eTN0I.D8C#f/J#>WHR<F<TBa_&a;_(/=-ARNE)EF>IG+J><fW]8X?5ZV7Fg
=MV2[g->^gde<DH2FB(WU<CZ\@I7VMS:@f<8c+GMe8AC^])M,U?O8bRGWT>N@5M4
fDG2Z#K/M6;GBXV?c=^H=+&b=/Z/:[=G&F0B/++Td-fX<SJfb5^IBG[_OCaI(]_K
S(Z3&FEd)ZB]gKI:&5M)W4&=Q-]b5UA?&fVMEe<I;2B]c?0KOfP:VBN5M.506J0F
V_BJfa:N33T4[0ITQ9;c](;Y(b9WJ1PK-G0@@#QCG1;aVW[Rg9.#8aGE^MCP5=/)
cb^G-aIc:U[B]LCd?Y.U0@L4IA<6A9cg#CO/6KV++J43><J^TT^J;#VI+U<1(X.;
>\XbQf>eg4#LXA^-^c<JOA3</H<^YdTC]_=50E;JFXaUZ#XC>8S]&5CG0H\?-E-<
1/\[?8F7]L5Z_[a/LG\-D-LZSU;MYB2ZE-[@HPDEA:RLV<Eb-W-#J:KJaN\N^-JN
&G_FBI?FBR1+YFW92\Jg\JDAJ^-/YF>K/g#WRJ-g2>;gb]V^;-4XU/_bCDQGPNVY
77).ETR/H70&D425\0<,LL2=_GP81YJ6I_?AUCcSMNgI-^@;D96U=g/FP_5Z1>4E
Z/#I4dYZaS.._V@Ba1?L\J2=6$
`endprotected
endmodule