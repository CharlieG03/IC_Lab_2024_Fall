// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"
`define PATNUM 100
`define SEED 8721
`define CYCLE_TIME 9
`define DEBUG 0

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
H#@O66eE-5D@EMJ<Sg&>6.Ra0Me)35_ZTX90PDAd;@BLDL_Z)UbW4)&7#S)8C&.b
/-088T_=aQ^R96S^a2,_e@N;F72@P7I-;F+RCMLUXBV7B5/6LR6d?L)+_9a:(X4:
QAQfb[T[&dZ>,eA\7OX:S-E<3T\ZX,^ESdEPZ(64PdPKO?MG^WX)-JYVDIUVO@8f
QfCWM4.ZBF6c)DO](<aX8M9FI\-H9=2H,Mb_&cJ_D^C]4fe>LR[DC_N>)?Jc-8P6
R5bD_.3_@AFd/B7[HKf7d>F#G_@_-7^?:NCM[g25]AL8.]LCUYb6G6;W+d>4ZMbL
T?0J><V8KM73bOBH.30\N=.G24Z9-]@T&R8ET+5B@VJ0(6LK+gE0YP8N539b=\T-
eI;W5-T?3BN8VeCRYgV_=\=V?BWHI;2CI71=]1;N)[#X@EHGGQXM_\VBdUO@TQ.>
bPGG1LFK_V#dPC.Ug=0UU_K8+bCgQbM26Q#LQU0GLe@MGLW+/I>L_-DKL?QL;ODS
9HQ?X[b7gPB,A9Y3?B[;^26?Eb,5=@X=7\059N2,Q92R;+JJ?6HPgff[,L^<f2WY
1I3+\WZ]>dS->CM9_U1,_DZ>/=6;V]f=L<ZNZ4/NNV\fUEVU#.><,E:g->1T=3[d
,L-XO^&]>KE4XVcVC=T_O73G[A\9^b;e(W0USM;9>9Rc@>DNM0]]A.>,&bHWXZ28
><\KN9,I\);+Ya@>CdNe^9;c5Q8:,F_I[?TY<F_1V:VD5?C:a,a=_@?HG[=&FH^^
Q)eaXTYJMg3.JbF[0)/>.b,e9:]=T\_d,FD46UF(95H29NOVQTU?b8]-=3[d/(X(
5.I64Wdg.(;:WL[S6+^AZUDYWN;O0/A\[&24d?:<2cIf@@#E)TSZNJISH0?O88=Y
HDV[.:LP(5cBfT\1&,=Gg-SOXDKAOd/VR./I>74^/XB&CEZ:ZHeM)1K:.LHCFONe
]Z-,PgaN;Z1f/L4GG693.74CFXe=>[V4a\OZ0Pg>eYD90SEgFg4=PA^?.YOF78D?
CEDW1VEKXL<O2=8dH8VIg1H\]b-CWGaMQBP-N9fCD9ab4T8NbCg[+P&V3P-P9/16
-ESRU8CA)H-Y5[8bc=UP5Kb@.](6H?Qg+]c0:D3d=2:(XXa?:+#H^VR#2+6@3K5Y
Ab\/<D=0KgMGOKLY?D=QXV6AaS#;\[1]W:O5T4&\;D:[:?/-A<@8[&UVV)RY1;H/
LMH[fNU+.)&_VS->.CWc9&N&;F>b5]IYC1-<(.LV/I/\e;?H)@+L-IV_5)DO:WM5
2-#JCEUH+4=72OWdDcYCg/S9,L9XgOI\eQT\&@BKLLVNS75V+A=]OHP-X[&XW7dW
/:HN-P:X\/GVYaJ5/DS+7Ob#EI\gV5[U0e=gVb<LR#>=,Hg;16aHI33>MXFA)\W.
Tf6/KC8cG2_XT3F]G4F7:,Eg,,4?QV/7TR.b8]Xf(B2MNT?4J^fM6SBE5W#2c4)a
6(4;EF-+_).-a.DXHD#d3EdXMdOZZ+WPeRTNHFc8A_:S34M9]acXXV[(5A__.,0?
2U@#344Z7?c?TQ;/)\INT<+Gd@-eADfCNG]\?&PZ[L>T8HbRP/2LZ\\,2@WZ4fR#
2Gg2-F-XNd/M^aWAUB5LJcK)T6GY7K96Z<-)HdZY+DA7<<8VgEeeUI1.Q4+N5,LJ
=O(b185U&9#;@O;[#R5CJO(BQ=d3>Q<(W6&->DaPJXT>1W9)HAJ0\0979EGGN=60
<8XA6b(\)+?LgF8G9ZG[H5b9G[ObK-f8;OZN5P3J:^ACXMV.gg.AXMQ\bZ0X@R.G
6:\ZPDH^.a27d=ZSS#U6B2RDMW5^MPb\gOAD]KJ_]3?^IWc6G77<<J(29>7c+[OU
/D]/S(;-Se)Za7HY@:AQ/#(5+Z[-F89;^AfWU^DX=gZ;N;WX43)N@#9QRWHVSCS)
W7OF_6<bM)0._I7\OTTE4/:[8=CDV6@I1=^3UT@+J#a^2Y[.N]DK[d07e-KW-[LG
P#gH#KF-WK1])S)DGXKB;a8E?)<RDY<b;+_0dF0+#OeCE#PCCLf3RXV?BMd)3NL8
Pb-eIM+6Jaf6S-c7eQOB;,T7fcPS&A<1gbPf1>U-4Ue1VY]6QBffId)J/Kc;K&,6
+;CRP2fBS,_,WP/B&Q(@C,=@RFYX]@R/>\(P.8E3+1PV2++[e^bV3M7NZgR0agMe
R8O6:5dYFK8c]bD6X+d.>4(]5]=>)KaQONc6^-7GL+.35+-=8c,NJ2\07gHZN0Ng
A[IG>(W_AXcC5@Y=@)Ig2PKDQU&VZKYI0U6O=gML@H:G=NMf78C(&)K\6ZS^LWcd
=94]gg[H&PRT6B>BJQEXP/XScfBOVE5C1Z>45XL+H]_8a&f@2Fa@+^[H/TT@DR.5
3#LHZ=Kf.Oa_Q.e9N?PI^)+M^Of5SOg@#?MD&IgR+D24QLVfGc,.=F)e_#Bd-PV^
Yf/eD<0eQ1K[0W(797?a9KPOYBZ)]:))@&>;B__+ETb(PLHM8/c<GZ>\C](<(@K7
O]\fFQbS7C=85P[ZBTAffa.^NB_1PdE^X&55,gWFYQMQ=<VB+D&<8>X5c.eMU@<b
4&VL;Bf041+U[,#CT[+Z,4QY>.W6dW)]VZV\J5N85.C\JF;]_(.H7:WDNH4-)LaU
WD#gQ7W_eWf3?8PJT/6d1[,YQg;UJ9MS]-+Z,FfO6aAa&[B](R4A?U>KTZ3<L/:-
X_L9?S:Gg(Aca\e1.=?[QPeOX\ZGfOZg-[:);RLNfVP6-R,e=0=JU^]daF>^a;7\
7SUX?96PgU5dH0dcIBQ:U2A@W/8:,-C#9G^NEY<gLc4Z9,R74VU=>6H^&)17WX6N
21M^EJMdL\R0,]a,B.+6gXcEN/,^K9RPWMW>FeF4C@(GHTCc&;@V)(TEgJa(3#aM
EIHb&aLdW4K2R_[=;g+._>=SC:LRcgU@<afOLc](aE)L+H.H#RDfX.eXVQY6ACJ3
;c_d_Z(9O^4666U,:-2gUQce++OHceU;P65NL.0d0UUS&WIUSb;LYW@VT/9\F=\X
,CG^S\4?d4LO+AL&\097UJP.AXc4Le3(J:7OE4<501W-26,3+XOY7)1Y@_7?])dH
Q(5XK88KZg,595\^4bJL+b[)GJ_YA6I2JG0HRI5JXL\F6bWXI4/Z^V&>:EW3/;Sg
6O8>4WXJ3.,[ZO&R&H43YCGWL(<\ScN42Fd>\JSULWeDL.PR6NVMUT+,VS6SKbMT
>7M4=<d<B@GU1XY-f@[>L=?A9_PadKZZ23+GVHeI5AMDS^K;0<QHf6?5e3KXN38G
CEKbV.Z^+KERfR4?O:,K<7dDN5U0QbC9VeL];Tg-UG\Ug]4O,8QG;#\[Y]E@?07U
1MM\cP=Hg<H)ID9V0(0d@WQf0/J4M;CA:O[)=]Q)aOSafC_4dVE(>Zb-F:?:-R/V
9DJT724GeG3)[-WEAXa5ZVZ=,WAG/d^ce8=gIV/d/,)LRA;J)X<(\\OY_cOCM<e^
GdA2O3QRT+X7^76J#f2T8DOKQ]VdV+D.(:>#dgM&<:U:&;.\MA_Dag1Oc>JC;HNV
3LD?>V=8G7S^)U^S]8-59JU)/g_&+^P)M]MFY-SA/BYdg\AdLLFKa9De8]=2.IMV
fP^=JN\LKeZ[f,@4W9\C9\0,)A=#/Df0(/NO?=X3\Oe4eB[d>4?T>fF\Wc89&4BC
;):WWUUAM5K=-cAJJ7Nd(#&YP51d4dg#?=GU^&E./=VYgYQEHR59,Ed]&8ffG#ID
CS1Yg41ZcR#2FeXN5K9R\L8g/IffgS@CW)UVe=NWW7TGdBMJW4#3f^4)^?3Z1ZOV
aVSe)YYf[>a5O3V/U((2I,+D??&bORKU&YGe2WX[&+QVU[>aGE,=9LYE@1e9eQN>
WbYJ20b.1RgTJ)8d;>b0J\Q[SMgN\PUD5-2-&MA6Z1&RG@BM]\Q;GbfFO,FO5@J0
.V8dUOJE)<d9KcbO)P2SfOIVL9K]E[:<XS(015DGO2LK[I08V=-\NF<KI&D]GNA5
=I5Q/\1);THHVbS4;]GUFb#/IA3UK@JJA9_YFB-QQ^EZW]CM3Q(M56B:<Q2<K#E9
fg?M@DTA9)5POaLC[5/SZc1^(:Z9:B_TFA1&6BR2I,/F,X+EDZbU]]fRBE>K_g?C
,EF/P0J44_9HAA90F6f?#^XOdR._E.e5OZgO<WFY(SXP\X-.EIIQUP6C]/3f>;aK
9Q6:QT#/:E_g@MFFf^GNefLUdI=YR,MS8J\/eJ>UL??F,A^b-J;;F-8NAN,C0SLH
_fW8.Y-69@6JFE+4BDf<>b7M.;-#<C7.HaKQ<TNW>67cf[.\4S<g-1R2b3A2M>+J
]GP4&JFM;J53=)+3TSWgA8M=N\c@O+E9LIEX;D)FUfZ/>6d.BB3_A,]Dc-[(Y?.Y
@.WT^K:L.3AWgT24NB?eeCCb@?b/9@b5OV\:c+aEda.NE9HRb6@M,G@BTH,/&1)@
CE=&VFB3\I<JQ80I2U0:_(6e):g4a&R(HV7Y>[A(P05F4O;GLYBF#:F^XgX-7\EI
)73f4/0/\.@b90QYWgW4?A06]LC7e>[ED0F:bIZ8[A?JWH.cG-[5XDM)&B=CH^EM
F0QP9gdf,PUg&Hg1Z^/-.Td@^9]S]U1:^L-?Yg42]\KC72L:UNN&/Z]a:S1O=(P8
;<F2]<ZcCT9#CP</Sc>X:JL:+A.U)D]ddT1B3/aB[I/a=0R_P]H:GFIXE(WC3F^2
f/2A9Q@ODe2QEH(NZIRV9@J5:ZW_GHB#Bca\E3a)[ac\FUER#S33+,eC&GMHSLRF
IXE&XDCJ8GN&S,E+^gG6RB6_9ZH6UF;ad7M,KUAEE8.YP?-S]V2\I3eUfe;@Xa?F
P2O:d0A.I(0aMP[LfVOK3Yf[g928KQ&(R->AXN]D0#UV</eI9).Og1PE)7_#+EdS
b2-4[>E.7EFF>RU6F3/D(ZT].5RQ,8<30_c@3>A4^X>Y>F&L<2A6G#4#/)XQ?7MZ
WL6A;/Dgc;0MH,<-@UeY<_5WbQKD7.dH(?YU#=:.;+F6^DgJHPQQU5&I)+]N+KU(
;Va=[JY/)(,X+[2?0X+4LZgK9PfUW_DV+E6b(4EN?cA[QeYF.=33:SQ0a>/&)HI#
KZ259[Q6N0-K]7a2d-S+A.9Lg.;?dD3O:/)F11D\,+ffHV>=ZK()@&Y_<=2OgTK>
C]A>a)7+Z;DD9]LO9DcM?Q<;(8]&4.(H)W]KfQD91bZFS:C:W^KbSP-WHL8_0[#C
5^d??VYO<2P]CR;8Me:a?CFVT<&WU>GM.__P>;gQN446L.Y?/B2S4+C\5=Vf6dE)
>E1)I(f..+&XSZ^b=N8aaORe8?_F0:+e5]U5a\F)K6;CDAaEP;[ML@D&WS;c1D(?
CJ5.2>N3(OC@-7Q8AG]?D&_8g(]4EKe+ccEK6@3RdA1E[R[B=R9T\/^.U[ZHe9J_
[(]#R4WP-A]X^./YM:3O8&:TC1+Y4CEb/YVD&G2S2dT<+J@cfFV[.[N)-/,]cc9U
4KDW9HUONfSPVOH9,QP3)<EYEWg5C_39dbF0RJA#Q>T-acN_7AVEC:aL6edS5AQ(
a<V929I8OUV#F\1,,+-@A3^XgAU[c+/EV)fB&CdACV&AV_QG59d84ZYR+>]G4&SH
EcW@D\6gL\5Oad&>O=2?25GSJR(&/?^WN]I=10M);8<C-&3KLDWT>T1JQ3]J4d0S
YaI4Sdc[(f<)OB?MCG?-._eCLQ#A.UN?b1++d.J^-Jg>QVWLKf_6#N:/_&R1g&@X
a;@W-BRe_72e_P8bf3H)gRRA2/MP\eZ]TKBY6T2e.4\YVB>2OY>agE;0V2Z/DHa(
3QgX/GZXY8\]bSZC,2G=EW1LQ=Y8^Q\L=JfJgJ>b.6f02A6>X#AN^.@\\V?U;-.I
P6P3):gZgK>JVR0(:S9@geaI.B4_W>[cQF.9+Z7QI5TG2^=GVAUAB(fV26NB_+X2
;FBggG7DMb+0O[U>2HRG1[:&O/HLC9K+_eGJOaCWUVfUFb/GB7U/PYNH4MI2)0&8
4g0C8:edg[ZH<f^K5g18W=1fHB(5<B1GWaCF@?E2,G4aR]<2(7:X:bVC(WJ^f-7O
0I42agf0@><b[B_8>Z<:8I33e]Ea;Xb&4MJKO4A.f(:Y=)8,R__SeYA@;c6-U]cD
\#=+Z&g-C=0N<24#GC8O(0OOaQ\6262Q4\:6H8<^<1QY41PG-&I-^@:-#W#8RgRN
5EeBUDUOM-@dgbKSU5e3XRH:R;S3Fd_0O2^?&R>]FSUOK5PSEC1^a@/V5(2CZf+,
J@bGE.BM?4<JGYWTD0K/@Y.POS[fc?\D;]],EX6Z[4Fe9PE4:/gS\5&ZfS^@7/J4
RFU+Kb3cWSaI0QZE-W_N&C\:g>K<(;I29U@YX()UFT3HMQYDWV+TgUCKKLF8Q2M9
#X\d36:Ia_d^E4PJ];151TdC/]Db2?0=f)9J&PV7YO=;PG?[3d^8,a2#ZMdgA?TS
50/gWNNK>:QPO0&TN-b,[<BcA\_g8+#g1/),MVW5G,:gD(;Q;<b=;ff01A:MV4Dc
I2GgR_d5(7ACNA254@,LM-T+gZ,fg>3.+0(F<?a:SH<0Z0TC3#1CPVMQU\30NO?_
409S)U:\WP00J(L4STWM//aPG4gDL,N+WC9dOEAQE0=d4,;I&AA[KIJ/F90UK/#M
_UU(b7be/M2[?PaCROba+I]aW1[fZR0G9+c(B@+dT-DL:-N:;Z?583XUF#:/PKMA
)[66:a^Q-0bf4T9C._33C(W#/V9J-S-TBE3#3a1PafJX6GKe5P,Q58F^[COG4;V1
7MM;egB4J=-#I8d5dBK8J+<)HYg32XV;@M=:D6+35M0DF3[@PdFdR-CD=I98bX+]
MX?BXTZ\RgBBW+PfCJN\P&RO^/LFQSB4FWdT#N@=+V#)UZH-C@S/<@[^BY?+T9[8
Y?2^#XM5V=3^fKXGQ(HL^EW?e9&30cPSVV-0DO0EDF]=\-ME,W3G/(b6B&HN_T;M
\1g>e7XSP_EV9&WA8>[D4>-WdX7RCBG4;fJ;cfWd3BPTJe8?f9_@cW)XW[5S_2)f
@#JTR]9KBLI\4aDd_UB\_d0ggJB68?OaK1K&2f>KM1a98bMPFBJ6NV->a0+CGZgD
L7PQ/ME37H69_1_P@,3bI2IT=V:D^.?_U9KA9YIU>K4W^/FR&A9J@QZZ8Y&&cY^f
=/+RIK7@,f1WP]RZ])P?\B7+U0&Fc\0;_:R625QcO=VU;&#D;)4CKQ40EB0-Cb\T
Y_^>DN^dXcWPfCFSdWd_F:L2Ag[HfPZ]CYM25ZEA53)@EZfT=Zb_-&@ebP\M^58g
_&(c_:,U=-22F7WBM,X[W^ObJc2c_#MB3#.X0<F3.SKE^1RZH;fT:Q3VMN5-AF6=
/(/KfH<@C\4#bHf<CK@T9NL#T-6>cQMN^_NH&-D_Z1:V:Kb]IG8RI@--M52BS[f^
UW^#]D4:bT6]J<b);\XI1M;GQdOc6<TC0Wc^-&VT.bY,(N^61K\<d9R3JAYZ&<_c
4HZ,gR&WKA:2:)LV0N\26F<(N\b]2C;GXT6Beb/2=H@WC&1B2fe^,LB/DMMaDOE<
?Aa(I1F[(ZZ2B4[JW^W4?.H#.FfXWZ)deU\87(:C?@A9H7V:]@6cOUU(bDGAfYT1
\,Yb54(@OD11(FMJ,?+,:_/9.H&YZQ7VBN\1\8Sc2RJ\Y3J^:/P=cY@4-5YcY]TF
./aZ&W.bT\/KLg56(MU=1W\d.IQ.]g-I4]/E[(,-PROb,V(+_NBQA06.cV_QWeO5
AAU.CfA=[1.ZGMDZA8K_J&E=Y0VLU8@_WZPfHT?3_409X.T+]5@WI64fdS>Ga3L3
f6&Y4?SXIZcSeP(gc[T(LF>:_J\(V;IFBTIU.#XMP3OUeX3K61<E^HPeIMU;1;7M
^)HP;_PPOM7.&3;2gW99(R+;;D=;M&TMEW+@;.[NeXUE[)F_J52,C;?Se,;aFBD-
5^f[>Ub<Y18TV))f1a6V9;b\RbV&a[UHg;A6P\]CWe+CHZY<WY<HQO44?P8+GHK5
-&S(-CZ-W4<e;Zefe+>(OL/CYaS1TY_\@7cX?W>.?KU\0_<-I;=?QBNe6ED9(d;)
;)Z4HUC3);TMSNT_1GK+FGHPO?>;YG<0L^W=Y?.W,d;-V,M\cacRb^R92POG;_LO
^W21Q6@)PfR?Y#ZJL--e#Q]51NQcX.2gN=?4A:RdAYD2QcS)<,14A9.PJX)FP(/V
T9C>TZCBWVHJD;d@LUdZdGCeRQ?cH;2PF5;I+K@Z;GQX.;UE[ZdJ^f_Bf_7B]ebF
W0f\1L?[[\fP+8+9dR>)7F0X5H;/IZ81(JF4NS,X4bK44BBf><fc=A@/b1)D4Z&9
5L]1eC;].V6=:f&[E4f8NB<bIVDBAYLQ\TVb^RI^ZF9\[88ZH^UX\[8RWgLIF&4-
7]HN&b1G)^>CJ\:39OVc/_CE_a=@754Lgf,Ob3+7]aD((g;RVc>D2N;^G?4H^G1C
D<_]cc6<?+S2H-<LHXPKR+6C>671W;NR0?0G&8#]HR=7da[:ARaa<c@7?S;-:D2+
aHW.0DLfVER,dT7A8@fcO<>GM#aGI2EBd=:ZI_]K65V/_RL?)eb:YJ(_-)Zc#V2E
d[XU9/ED@e6Y-S8D)JRR&B/?D-aD?XLA?GSa2DJAcR4&e@P]]W&+-50&>[8SQL#-
;.?.Q,7aNZ\LY]548FD@[(bedBM9/;[1IE^T.Z)/N(L:_7ec+b0&K,Y/D2ZI]<f9
4A->_J4WVXR.9&/[c4)KH&]]-:<P\YG5?a7;L^ZZUK/3T=QJL5Kg/LRe<4CBI_BU
B&9.=cOe?\M2ELU@@7-;0YO_N)BGJ7:-4??gbGW>#(=M.D=Vf2;)/B/&BWI(Z&<.
>8cY;bARa,b;<L(#DWeNBL)W0P;cO-C+?L#OJV^4PCA[-e2HA4B]6M_K:&+AUT],
8I4RfU@)>KPP2YNPWYHc]J-0@CHJeAM^1_6C7<e;K<c6Ze4#KARcO6NNA=5Q,:[_
+AI]R=GU55e;+S9)/#JWXE>?#T_9b;gTXI<:^_T7MA,]+4&>)&)#7JEWA1e9(VO7
E1dgFD<8&&FP;NeO9VVEPR2+b2VM359DXWd&d:(>D6;=PcTMZ()JLU1dS</#UHg0
VJM(;Z0_eTS?1]#5T4W.V;)A=ZW#L.4L>^3\5<]Z</g,e?V7-7,ZOW/7,:g,0=/0
AT4[0fg/ZZ?@N_[_8-V=[dDUDg]a^+KKBAXP&#7A@fS:ZSXd,,<V]0AWRW&<2g.2
Vg6#M@1,9)dXHC:eT==Y+&C31VZD>9e3O^YM&S4dd0(\>YV[[UQ?eg[H8GD.a[UX
AX328cFS=eRNZ-VV7((])5,afI_@UGG=+1;:Eb.7Qfb?6_IW6NPH)+=(W873C?8Q
?@_5g);>U#RZFdfV9S-&EMO@H:QNQ(bcU\>;2:K0cN7A+9<+BD8()A(>W@)I9?4_
>BNNC<M+-c>M./2d71>.:XBXf]]Y70XZ5,c+gcN?PMAU14M\UBU>H9APWYIX.^VQ
Z[<aUC/7M82J6U;W=dPK)8VR5PXG^f>UR&2M0&\fW74S44GR[WC48<CVCWI-]#MR
KSe9RX.S/GAL/>bG_KDYbgL+6A)B<OA+f.Y#K:_McN<ZL0B,g/D6D5TEVEaT\^f3
G2d1C:Be,,AP@2_5R(>eETdb2fUP_=A^(@-+F8R3T<&M9aWfe/D9-/^3/A=FIH4]
)OC09_OE4XX>eL(R]+A5^^V??OWR0c]b^Oa[9>]0WS0ARQ58Sg/OUL]VKD<fEFge
A.V+[><@8:,(4\A5(RF^\XNSB=(bFP0=,N=GGS?=,8IV[A_S>JLUb6bT;Nc<JVP;
RVX)L9PZ-Ue5ZGN08V+9?FCXE^NRJ\]14:(8UI_,BSGR9H3:&O.JYXJ5=&Q5D8F>
<<@DJIU\cXV@73daL^\HAe>OcPgfU>&S<WY>=TS0;J)T/M-;,VBN=gM2gd0N)fTd
T8,X]4\UP_)EX=D>F2Y2f\2gKcNX/8(MFWA]SSJQOba?4^9W(5EJ4((a4YL6EbA[
GL4\Z(Y.;UA38J3^FI#U,Gd=#O-5R:c@=U_LcLZg[G]a&O3J\:=H1#\1,DJ6I@QW
]Kf+/K_W+LB?NeO3K-92a.WU]PHK&7eLe0WDd4bPZ[J]5eFg\[FI/Y0D5f?Rg.F]
6B@/EVMK.]2ec/9XS]0Wf>)I-/?W9FP-3WMG44_5MP>G=IO+H\E85b[C@Yf))239
-;^PB[)^VA2L5gR^8P#7N+2V2YW6KbVYaHd[UARO;aHU4bR+)TM?4^.B[aXS@DaH
1Idd:9M6?F1I_8-VJ\:&+eS)-U/G:0UUI=+MRDZT;Q4bV,)H08:YAMH:ABEU+TUA
ER^K-//>bE)-^Q<PP6;_\_QYb36e2UERfb<ND\N7ZD0^fb6WIO91]ecL;Fc6&=YR
^1[3+YP>LDLMTeC5@HCVP0.5_a<2#@fIgUCL4T92I7_HKRNXHSC#^(\H]TeGEW<a
,Q_YB2YNX<W59WVVBBcf0]9;,YZ=X@WGN;MSeWP^1@@LXafaQ>b6AB.[\ddU<LW9
U1)2>Y46529CG+(CQ;XMdBQT3fX?VP<71-Y(Y=4e7:+eccJ9-&E4TK#PPc)F38gF
[_Ld)NS(XO5Xf(G)K/_R?gS9OHA38?K64?XG[\2]//,FOTUB+V.UJcd[12[/YD#H
CO:@K7[dBUKb2NHT-:,K+aEaOW@V/=DOCCL6(RZ_QSU[)-:_b33)SZ9/Vc7>B9LC
V_SeM+&Y>P#Lf3WRPGe+gL\.a7afW7O11U-/FN_1?X^JS6NUJ:D5</29E-]TcTC4
WV#TG4P6)O,93WD1V6I7--;GN/,aE7?cP?E(Wd[7WO??6.[.-3GWSYXTR<DKEg#>
CK)b@AWWgW)eHO>7B)J_Q\IN3PObEV.Fg#B]K(;^:D5_[eb:6?R\/^ZfQITJE7^>
)GOF;TM;[OUYHa9_E[]:J56YcaIY989SMF[35R233?J>E0ffcE;J]8-aE<,#)(03
T_N>OI.T7eWRWeQdO;B2\-BR4@111+VcXLHX18I8NU&(DHY/0a>P6@R;OZafe<0Z
LB=L1;E9/,IRB&05VX\5V3-#VW</4Gg78,52<6c#_R,M22PG=?S4#61&=SM?YE54
]4L12],,SQVbGOPKg4)7ec8EAA27^2ag?&1V4aK)@M_H17-JG&FKVSg8XWDA#R=/
\X^@HW;@RIMN>JH3+ReEJJcN->feVS<#CIYE_Q(N&RSG_EU4;3-PBA85(?La;6ae
ANg_T.-^RRZgJB]aA&b3;3OJbGNGaOQ.F+?6R/UK3Keebe@SM&&]aceQHJ,>L]TY
S=&aIBAY>MP2BNY-92_FT]MCRPBC1>I=9=]CE=&_AWNA@b?M;S]4X-GOVNAKcM^K
1<H:4HEc?HN/S/)C3<Qa?MGS;:&@;X8S&^O__G_6D20<GW#gI@^dZMaO-SQX=[TQ
J;CX8gK8ZO:F306,H>:,BONJL;H^f/0\;^W)f_VF1@7/4)<-60[PMFK<6YOdG,#?
??FWCPJB@aX?#.=R\IU@D/fa8^IFH.F03dD=+,1CX[I:7+7GB@,&dXZ9]GOF8U#&
-BZP<<M=U>PcB=K[=O:<=+,G\);<a9W3)]]AHfI\A^DNS3V,&MQ6cVOC:MWUbEN+
;LMC(ZI(8N&#5ILg#M;4V)HH/3QQ<H:UE&b8E@bWTd_)ZC/[NDHT-?/2>#&geV(d
.8E.g;>a[._/@)+-[I9Lb-,JdY8e]c#D,?FgfKS[BGQ[M4082B]0@Q^,NZOgZgN8
GOUBI.>2SYX_+6B+5Sf#J[CXK?db5(8RC<fAaASF7#<Rc&OLCR?UT<&b5^dY6b?_
B&2gX?^Z&eP+]71A8P][IAY6VB.2Q]d8.c@;>+;bK+>-Ka(+,FT]bS:H9S3EVK4>
+R,7I8EaEZ9JNTK#SYf/PZ=4RAHG^Z)&8b?@5fVSM5Q+CP#V;3CWf:+QeX@,=;NV
1VG<^\QQMR8+,X9&dB?F<UE8A(=\8PRdQR\&]72^-[I,;-Wg5=1g2U<a+B;06WP/
IcZ34&0X99b0Q/#gGcIQdOHF4<c&E9#85eD4R-5-S0):Ydfb7YfS[e5NCB3@@]dT
+]UIb#G7D,C<8@;RJDT[#^BZ0[V^[=3/#45_DX1ZY7MP\VFafST[e^@C0RWbEdUb
FJ,R>1@_06bT@XH,:=8/cB8+Y9+<@EMBHDMMJ(JQA?B.B(\VS95O\+ORD3e)G&XQ
d4?Y/C<CMKS0f/IGQRcFON8?B7(>XEOLZYX0KJ8L<0fY7=MGM0dZ+X=T>FH,HW7e
Z#FHREbe>B_5S0-OgRf:]F<BB_E@;?V2;YU[W6BLfW?5G=/NAN3AYH,]SF,9)ZK,
@gINPVZf^+\[7]T52=,]:-Y>[DM3df^-LZ??..)W5)KBGf#FgM90eA+Aa9/8K5E5
ddV)W(X^/Na,>aA)+\?IEL0PWb)f?RT>J?BJG\PR95]S[_;=GG/ZT#L3X;.,KD]E
LHAf5?:^YB(GB@b;0ecV@9]J)OE+-NU:2N61e\(;RDG4f8=>.?Mg-4)^bUBgS(#/
V3TXOD3eL&I54+@d[Q(DL>Q,H;HLH\FU+N0BL1R=A2c:I4?X/#_\;0cUe)4P0<bf
8+;J;VSO#.OZVPgC><CW8)?CbH@V,5Wgb@M/3OGg<\]\S2IUbaQ>&g?AI6+P:T:c
T?/Q-I/;\Y)&A/A(LH;88-8R2QHF;ZF>E@+f;S6H#H0ZDO8AV?LR/cC>76_/O3(8
-QPZPJ6^91_<#NW(;Q>e+PRbGBW6I@D&ANHdH5>80SJc2TW6.b)e,<BUac10<gc.
I?G>:JaeO5NBWRYde-<&g/gDBA2?_8NPNO@&9S]dA.EWJ=<.#<\.6d9d6E)dUT?>
K8aL.\=,?I=EY_aAbU4ZYN#HT#?9P^2II4=FZQ3>_^;R^^83[3B,.LB3ZP.9PW8<
FdF+0Y_5CbTL?B6WU\QKV):;E)HHEfPTf#5TeP[g>XH:T[0>G-\9CRHc+[^T]FD<
Za+Yc&e^Z[bK#=6T[b4dI](>^Mg]-I1_ZJ#>[)5L\B0e]cY1]_?DA/,8GZFL#25)
b>2)+(J5ORPW1DE3e__Fd=FOCf6[D;EUe0-U+.XTS2g+(N5.?.36dGGLb@HX[K5)
U@Y82^7?\8f,LG;E.BY?BL=,T=)3Z\-,:379[JZ0)M?32)/CPP5926P^&>JX_&U1
8>RNZV#C20[6abWUfPJGC5^K96+cK2XZ\57:HASf)a79<?;cBV,/+<bU(]6\7LZ\
E_Q8Y\^YFMET-bL?-XP_2Of)&6]6FUMX9>CIN_XgOSMN7=IBAGB9MW[<7BSaA#@R
,&2,b@19a[72(aI<Ac];Mfg^KHYeRNW2J?>RT4#(ZTT8(9BdU&52=\,f^ebC&[QA
VeNdIZQ6f)89YH7#K@?3?9XE]+8ZAfB@?WFd&SQ7+2I[I^V[cNaO@32^2cLY17E)
;]1c,K.(e79RJU;?X+=\HPE?,EY;PO=9Y_D]_FT:+OcB_gH43U72+S(1^==V@d88
c;(2eFAdLA6U0P6V__YcK)M9OQ]=N9,6P98),VD.LPC8Y_O?+K#Z]^e8F71V)86S
)Xa#A.f<]G)MNbR/Cd6GMfW9G,G-f\H\JeJ>.6HO0cB3M30d<D-,Ne@.bX(+:/V\
T01X,BD#+H-g@]2G\;G9PA\VDM75XVFFP#6N(]QW]E53O2fRV9^0[AA4HeT[K<T&
30#LK0Y1,?TU;4:L[5YK(_^U&?7:/3R@&8Vc7\gX+:PQXO]\GZ8898,?BOa12?e[
&/OW]9LDf>Ld,B2=d@N;G#)\fH:AK[[MK.&9V3-ML:QeYTeX<(::DXUeD0b\@gV+
>R>e7I/X7;b:@L-_]LR6+V:_02/[G&5[2VS4+TXI.LP?Rd0.C^dBS.ZM)+b5#P6Q
\[-d&M;N/PSNQJ>>Mga6+-\(EN,9-f,43,+@e#-1&@4?(Vb=2.9;eQ8Gc)d_8,RU
MCN)^:QE75JGUfSSADKZaeMQ.GbX]LKQ^D1V(fd?eBEG[YO7U#.0<;.FQY(=V=D[
MID)G1L]08[Q48cQEZ@fF@WQ[Q/(5-U[Q/4E(T,O-Aa)-CT-f@6[,aC^2H:-/e]R
+E.g2M>AL#;)N^AA25eK2-^HVO&F\[#T;QGJ(Z)WWJIAL33W(cYN\U:KW/aFCY?H
5@D<cJR^Y3_,QY36=8.c7bWK6[=/5NK&fHQd-g2P=Ec)20]C8X,>5=eAd4+)SX7/
V>@?Pg7T0IL)TPT,g?UQ_CELY:_;ET@+VXXb7P45Hf20]gS?HLPN>1CU=;9.J0HT
;Xga4#0?,^f/8f^S.5Rc[Z47e5C3-2a,2&2X;9G=YHLKV>P:(Q13faEK2T]Uc17V
eP&T3<;U_I)c#OK3b@g#e48eHE@/94S:E;W#F.C&UK1>^5F&fZZ>QWQXS>RE0Hc)
SX@_eQ)ZW?FWA/1DeZaOF@f=4@QK3g=G4S[S8JN#df+SG8d\AYcJM85YF0OZ4d5/
1PE7d#?>1)@,>Q5[-94HJ:7/@5bFf+YU/P7ZD5a)3.1Lc79[TAVE@YYI&XLZ\6?3
Z2()3<]@S]bL3N>Gf.6-Z]NRETfML2QW)MAd5M6cZKX5TO/d[J@0aVZId^MW#+#T
+H9Ke7AabRVCI-bR9A2#-O4QR5M:L&C<=A31:]1[[7I4f>.d@:eO.a8e22Q_e+B^
cGL>ZN/^&_7XQ^+2-Af-5d\cC,<Xcg63e35FF&G+./&f]3U@AOVVB:=2DbI>O0WJ
(R;@64-^D:Y=OO-8Z^3KE_gGWZXK3IT]EFXC,,K41=#abaDJTc.a&,6J[+LaWTaS
cV>/1[6W39CRDaE]L2PSa=G#@df2P@-.gZQ6_R>;bT;VIT[,_4EVM,3J2(QI:&OA
_FT2A_HRe<)W[[1^IGeeJ26)U_FceT4S<&1eK\Ed-eSA0I.F&>;RPgL,#)F/[VDJ
\AB_6QF9WY]4LJ#_Ge5@DA6(#^8bJ)a:QDMd7=CKR2&U-)9Y1.0&0PM=3S>VX2M&
/Q&7JY]9&EM?A@7J+?2(#8[+U<H&H)<?fH1E;S2.2@?.1_UV(K<bb.N/NAE+A(EG
Y/?34<FF4K)8AMf,0Ae&]EGW_IUg9-H,A:;T10.9364NTYU;+W>=[948N;?A+>^X
A#-9+b6BA)8SHLLREZ?T&&3E+ILU53cVW+\H(aX#A##2DBEBfVd@]3VbPR=B&CQ5
JHD.2TCD9c,+,VcN>U2F+g-IEXFI;7_B(GJg#/UE)f_4JF45_40M1B.ST0bMDce#
02LHXB/;M-2:WCQ-FM2.B_T=.Ge5bF/[48W2,\/\1eg@RM[HNVDB54]]:^;TbK7f
L8a;Kb#\g9J?7JeNS@d12=/S-cQ=UFb_9IQI3;VK0(SA;WO=a(YHWf#2;X_ACE/?
C2U_)LN@Y0KaF,BN;4\J]4B-D2;Y@([OE<:c<S/\YQZH=>1H4@AR<(Q7D5PHc/[Y
+4Ff>K4#HZeWa.FI=H,dadS8=LRgW<L=QNTJbOZBMf:,e-\OVf,=_7JHG^6Dd]PO
VS))HR->dK7_JCC2[R8(e\c\EOOb276\/WfC].M4;NGO6/.d0=3)DfR&HS#BeQcQ
]9H3c60:eUN:,P&]=Ub&1P0bEI].b#@YCbQR_g>Q)gMJ^A7fD<_[_B#99H2@IL<]
>KRFF=b0?>NAL,@1:L,?+2fLL0e>>4P:RRIUJXS5EO7;CY/e)#fb>#XWbdAW4&A:
@HQG1ZVL&d;YPcKCXMH;Q+?V\Kb]e\-Yfc)^X:P:F^)DGR5bN2>ZdC=[0&6<>5e<
OAAbgQR#&5,YOc)JCSL83TN]&5))X;g7_NW2I7LGYT04H+L7GIX7MZ7O[[U5fCVI
,>de/^L9FG>D\L6c2X=cgUCQO+247SB[Y.PK1P_]^]B&XA@c70.7:-;27)PX(&KD
\d6O)5\\.9]bSSD3f+f0a_<->#[2S(W01L4^??=ca8)#5+.e9C@E(846+/B4e8C@
0<)_D4=[)0bI/aCWbZVJaCTF02b3Y4P(I/ADfH]@9\6?/:\W]@HZM4Ja0Q[1OF+L
Cd^fQPNK:e..FCe#CBC:BW=\RNeBf&.<Td_..S>QR8=f+^MY\FGYXCK4Y(\)NZTg
C=MV]KaSAeT#QE3HaLBe^,DFV0+ANBY(0XVDM]D/]CO8gg^0ABK6A]&UW4F&b:#J
ff-[J,WZQ_,3KW;]0A0A2=7V7V(Z2:SK@e6/cLaKW,2SLOTARU:K&d_e@B3Y)316
C9O1S891M@1JS8@Mc0-J.VTf(GFB-4E9B[RY@[d61?M.9;)4AIG.Eb&Hf(<=)Q]C
C:=eGS@58PIVH]&[>(U.fPMSNbVIQ;_6R9N/SbQ04FT-G,PTMO(.1Q+VBRL-YB6R
_?I9<&7=bZVUJ?-:IYW?ZK.(fY;6..WGD\C3TV72gdA24W15Xb;XQM8gP,SCfBa-
>e@A+K9VL,3[5K(dIN>,];9WZ_e8LHJ1:)R+-d@#R3[9W]@V,P-X)MFVD0O:0+^U
^3=R?(WSQ=gWKL/3JbIbC;,;P.RL-Ad.6P?2+RSdE#]==VfFIKM;?0U@V4+XZ0(<
7?64UGB:c0@_S,D&f2O?d8U2-ZC4<a.M0Vdb@C7YaQI\0Y,/F@NB5aXaS.K4@fFT
ZWNQMS]f3N][LCg2b6g-G-ER#6g][H1Z8VZ/0SQHGVKZID?8IJUfV9&+\)5]O:Gb
Z]b1PTV>Be0;RN2Z?d(B23U;H],ED6L2</R^X8(7LQIP:]2H/<SSZL,RL\00#1LX
QK_HaE-ag]2S=UZ-?C&dP>P9U6eE6IHR_RYS\_dHe_ZfFI64C4dIcI>M>?OI?C\.
PGb(<D(d\WfW5DJ0A[XJOLZQW=-\K+V4Q43fD,YOT>RbaWSI[6E_3[F@cY;cEV9@
@I7X?5AY0N&gSW?<;BE3_4&g#H?6b@E?JJggZ)..0>MNK,.Y_fWe/[(b6F\9O_/g
6G.[5D8UC9TKP>Y[6_?2_TU:M)de@\XD+PSXaF.K/ZWWPgcCc&:.?fM2<@IAKJS[
eT__/-@#;0_g:fLR3eWX?,E:JQSQ4fX79-[WO/7(8dNMJZ_URMa&Jc5<TGf@V75b
]S-/<\.SJf2.XI]:MU8SD)#G^\R::7AUHD&YUNQZ\)_\6e>SK9.N&J@,Y[f2b<YU
&K-(9P@DTAEK[bec]0PD_JK:,SeT25TEXLJ6AE+XRLZ1^K;I@^Zc0dFK.K7LG_S6
XP?Q5)d+)NUcP>a9-#Lf-Z45d,e)aKAJQGBJAPFfG:HXR5K0beaK:94OeI44IU;0
V8J6S5/4ZP>\;V9G3dYQF9D7#K)[<1=>Za[H13Z4N#S_H4-9NaRDEPaCOXXH>[7>
_HCRdVINKMWCV.ba>.UTMK]eQKeF2fLaD8Oa3K7fD-7\E,,F,P+ZcR5;-f1<\eWg
CBY;:YL[V7Hbe/Q?ZY)/UMDfdZQV]TQRP<O3I_Vfc]<+OdP7@Dcd9d6b1Ha,A[RS
d]BR&cYP;_W#=B?@97]KDZ90]1OZ]E@N8?@(^4]X#aCKD5&a[@BKb(P^VA6@D>-D
B=LE71/T,5^D;6TH7]I)AELbS,78^YcX)Gc0H#TR=:DXFVMZQQ8F/BRHZO_NaB3]
>[JMEUQ(YaJDGDG(X;21XWC-?QR7I82#CIR2&G;^DgON1;#[IFHAd.=6&Y<-@/=9
M9;<,_f9XQT1X?,YC+ScEV_5GOQNFX7V.+,O1./,;(c(e5SUP0IRPO<T8LW,f-HU
?UTV^=1U9_NLI<_d+_&Q[?<98]F2EdJI+=be<^W-916VSNI:,\03YEH.7HV>SZSN
ge@68<g7gC741_.1Fd;M(:P>bJ/a1P333M0.09:gLF0Uea^F+DF?78;a@@2XSLXg
C6,+AKW7YTN)??5VJaaJB3.TZb_IZ3Q/#g^3K2WAI2U1XJ08a^-0W17N=B>])O>[
_c@&5DJJea+>N#[E3]9,R?dTO]O5;,;]KAOO7ORD5JRND[(I6>6.OSb+DX7[g\ef
CR5X7d7:=80VTSF^C/CW3caD+c)UB-R#R=25eZ9dQSD[I8Xe3J9/f@[a@?\gLN^d
GAOEWZ<O@8[DTJ)#-2[_>WE+G(/QH/[gcO=1gY@EO[QQ\<J]eQ1^cA_@=],9AF33
>7d^\IT]4V/-A_^&??C_B73f[2_2DB_:KEH.)/Hd<SVKAL\V8?1=RW-@4U9?@bVZ
SHVYXZQ9eH//JIIO2X&Z#26?Qb6,KTL1-JW_c<T)BYSBIB-&.?+VH#N1EU6TH;F0
2P1]C7&#3bW)Mf^6W2=?YAGY.;,ZdR/=IYVIN=KeC?b[E12OfFTI929NDM^C<;13
AR,)F5I-<4CO@-d5ScH-G/Lgf>[)9+D-&W5bKZE&_)-^[5</:2]3UGR#VG3AI-@8
;?4Cf0CJTTA&c3W5MV)<8TJX,Y#-U^cX(<4D_4AT<805bYXP7W4I^3g4IVO@P1AS
(P2UAgBX:U0BKWDKb<Q13g]X_T-#+,NdE^LD4YBb46FR3C:X.cdTZ##\1K\E,g@C
@LT<MMf2Q7:@^FK@EdIFX@?dLJ=1@Z?-S>:@JYO?CUXL75fA\d(E(XG,c<0YQ7/B
PQ25<R\RaOZC7a.fR)?_V0X=#gM2bUPRX#]ZHDN@6Q06W-RO):c7^AYJ1/^F405H
EWW=PYKJ/B.XbV/9\.70#8.,[Ja)a)bK94CRKSKZC_b>JC\3-761C#\XWE_,C;&+
S+DT;AM_D0(T+gbA7&BO=W<2+YPILP@5cMPI\V&\3_g+@fNQ0K;Eb2NJNH:F/PdZ
_A8^S]Gde:4cQ/FE2)4M@<Q&-Tf?W?[R5gOY027A2S,YMBQZ<;228YNEKe^ERBdP
2AHK2-:1.?>=4U><9aGF23ed<HI17#EH[c2.4?>.I8A\=R,Tf[NBI9ObJ._P,-[=
SIgHLe_20_X(^:V0bAAHUMAXd\>NTbL(>-KF-A\Q,,B+UYU5HETTE@B2GAOJ0D-a
OS0.4QGc>J[GO_bLS[XW,X8P?7VOJT4GH@#MU9SCeKgL7I+7,,)-0I48ZXN+P4JS
a;3GW@VN??G1]6V4P9aXLJ_M-@Wc>A&Y./ge)/B^9ZPb0A):A2F@U+Wa\E+bY8V-
]\aTQLGAO1-[BO6-I9(W<3QZbM+2=8(9]AHSRdSTVcYVf9<X^Ac?:?8+RTSda>WK
)>X+].JJXFS,72?SU3IeO9AW##/O58OL\OR-;3#J=H/=dU<3KTK(db#CF^XWAdDD
/^P7<87R:D11,H+HaC@NK,/gVbO&+dbXV8aM2K&4@@TO))DcHUOZ<\6>Y4=4;LF7
UO41RUIMH]L1J6FW6/YFKT?NGKT=97g<6\WM6e)DFWPSaG^BdRHb:]7/Badf[JRY
TO=HXE2>,?,KL@YFbEV@/7CI9)?Q7J;GWCVR1+K#CGBUcC(G2e524?NAZ.0Xf9g0
2,JV4&Y([U[_Fd8\H,-.4gU^.aBU2(U^(=ES(eOVIcCcEe6I6;(Y9P7KU4DI.&7f
&S?aL&[RW3;F^RFV(09LMK9^,=_T;-1A2^^d_79\;\BW<3CT<\(M@[]81]c@[-?A
;-E[RBe#FHfKdR^I##X>g@L4;\dV)IHQE6=(b74,D2b3e,JNR8dDD[S/CbHMXT.5
)(@LWEW&24=WcXWO2?d3T9[P#;D#J=U\(IC2gRQ&J:-=(P;P4gg>&Jd;a)@IWRGB
):C42BMO_WK5U>a;=feIIOA/)(:GK(968A3(DP5-J5:Y[<T-+=GSB;XCYDULe.c)
[)975@gH)OMRQSe9(6H[QI71P^=OX8TZ4FL8T2^JX&Ff[AIY9ZK;7;.)DgI1d-Gg
DE73>O<f=)]:?+g=SVT4FIPL8Y@c3H[eZaTL6b.8(Ea>:MLdd,b,GP,dQS3@],QA
G@^TdG//XZ>3AXT1\B77^-?<QW0F8K@FI/;KE2PeA0]H?6&,4bNN1C[)XNAc)IZ#
3VM_Y]-N)B:_g74BDX]AIJV>a0E[:ITT@B5)Id\aVUbL\PO_VI;/NYeU.>=<]9B1
STQZ)9-U>T:^<3&76e,F@/f_FWQ/1^RY+OeB#A0S-OG=TK9/FR_+cMK4N9363&.b
&K/31>^LGeY+TGGZL3^&K/E:)##U532A<,e<KY@BNJX4aSbLb;++&Eg>P;dF:;Da
=Q4QgJK^\6,e7?+_,SG.C77:D<N>ZPQN)@B?PF&10A/cV>=PSF(1?PaJC/I=PP+S
b3&=+=NY[/;9O_?I2WPg5GCd&Q[c@PLHFad]Za,7c3M^;\<DaRd<UK++XeMVZPJA
#DAUf<<:SBPQ1f\/6^(5,R3?=(V_,BfWGX8FQOH;>UJ.S1W.DKafM>S:Sd0?:^S.
WB;B8&(7\gf[0WeQ?NL1UN@WNBWfES5FU[eUdEL-3QH,d-3F)@#.f5]#V^J],Wa#
;bR9de;b;P^Zf\4Y2+HV37A20d<2>9+cECJ[4.^af\HIT&8Y.GbNC,ML2&AYN5<T
SDDdFc(E9:G6Z2?U<Ed@)ReS+2YB7M;ZWG]=1\CYV[E(D)7BDgYZJQ/@])aV:ce3
-H>N(35MOABIP92Db++f\G.CbSDG8G=@-TL5KO78e3(654T+3/cN#9G^gV4bL(/+
?GJ1AW=_>6;/g5-<c7e7#MDU5-cGS-@8gbdV:(&P#AX+X(Eb)6B0C7\(N8Q37dSM
b;W_Vg8.LVSJ1Xe3Jef;gXYK10HKV\POQ4ba1:&^U1a#^7V)>4fbR-;8\:ge,S;]
Wb5cEAMSGa:L2[c>,;(gSNCDH2PYW.46/&9HIW6XdRdJNg#>1TA[.)@?F_gTP)1#
c/aF.CMWRS_9R(]AcK.^HdPU+NP@dHZSf&1Y\=+U>2-W+YFK:AL>d_<47A3RBR:b
VS5UWfG2.8):LX17?g6,]#I^2<6PXP+<.7I2PPIKL0;[5PA<9\>,c)/Obc\02I<(
0XML2HVH:&A[bH)?)+EH8:;1,,O;eTY44G5M3ccCdH>]^VH4+YQ]^E8IE78Td@?e
P_]IGX\R-VL&<\WIF3PB:b(#)XP>OC3^GP;86Q1#@Y@EU/CB^(fV)-3;ZP#cAEYf
#PIeA<6:>#-Q5&ae07\ZLRE\+?U1\Mf?&6V37N+LK<@8#;C8YB)#dSHKI8bFMS^#
OB5bEF+LD4WT?#BER9BQNCT5V<.H^?,BK)>:-JgE7+R9SF0Z#<T7FIdT)(K40J@#
,&@B;&UbE\+HIF<TGG0JPK>YC_;A@e]-4_a[9Z2Yfg7;;K2&b_&<Z>dK;0XB<gM(
-Kd8EcPBaeK4<(QaAf-T4M4b]]E4Q1TdURbIY=cA9.]?.+XB#(P,9;fJd&=TM-Y]
f8H4I-:ETgLO@.@G?77[Wfd00=YC0AR4=H:+E#E6M^#1;)T]A,7#;2gK?#N;&PEB
X9@^bbLN+3d3W)S<OH<EX+&@4GPMV=G=7Z1#6;+\9c8[AO5&(#]YHfIF_;D;PB-H
<JF\f2a:Mf17N;N-bV,;O,8?c5I06Q&P)W(:XMY+8,>?>Z(&+@RAZ)aCKU3+d8,3
\XFU3gZa+6eEZ31PDE1NV^-<L/5=OL5=aCTBY+&?eF#.,>.cW<=]<S.&c(Qg,>cJ
B,RJf:FE#fYPeC9QKZRBFOV,(O^PR5C\f\)NXO@AX./U[6/8GKQ0AD-B3&VKO]dL
-L-d4V5FVLQ8)5c-e&Bb+-UNcV)?.R8Zfb1IccR+ec:,1?@29;03Ng5A@>:#CEc+
#FC1J25La86-b@,](GTQ4+86NXJQ17&UOf\VY\L757[5XNfNZ#IYI0X3?UH7B^\a
>JHAD];E3[dAe=/,.X4b>\g8+X,P7C8_#DbIF:W.acL5Z:9^D#;e1F4+IZ2_0/2_
2N.,:9MM1<]4K3ad_6[3a,,adS?9(B7K_SVIBL8N[GLYXFJ.N/VbKfg@N?1d,;/_
1aT[(Ie8,.&dc?;D<Hc?UK_UK<;T3HafY1]D>J1[Q2H+f+H?FT=aEJ59e&]Q)4^N
O6Y2K<;CfW/7_H9MECN4<R\cAI7#a,W2J3bUJ2)6E6Y#3NcbZU<Q79],9/<1=+RK
N2CcZGKLH9R+&>=7LM\<@-7HG>c]23I3bJEB3_/A^(NOBf=)@5G_OL?JCMLALCdI
_LOEOVWf6b\5@gV/NI,T3VZ.LW7IDUE#>ZCE/^A^LMag-/XP^,d-b+fJ,2)>PI.F
W+0&F2\H^;BA5C/>-c9fIQ+@8FPQO8d@Z4Y)/<OO6APGX8g&a;F6SAXBX[VK\TLB
+E5Y]\FO0>I1<SFC(J_dK/RU\c7&]V0#de^[g&PP0V9>3J)I4/d?XU@F-bP[Z3?3
G?ddRUWUIG[&7P4]TSX0ZW2OB7]1I+O_^4ff)3MN,T<CZIQfa8I.Re)0aAKU>5UX
J&9M+1AT(gQcIf^Y[G^EEg@U\2S<I&&CDJ,f:If=dSF4fZ37U7+G2[9_.3I0aIJF
\IIa,@]8<^\H>I/=f]dSM-LK,AL/G3&Xe-9=.U;cE0E]C^U4B+@-7;f3#Z)9[AGJ
=(K;?PE::?KJWEA3B&58?[^V[gWD(g2ZOR@F[Y1dC@SK-AT-fT_NSO2]R8U^3HP6
ce\2U4\>LW_B#+gYJ\1>KQ\_<P,@2V<9&_7T-(=6IP,0T.5W0>YUI#9B_II&EQSM
d1aW\;-T@)=KOKf)TSR?^fY+-0YH&>W,I5E1)Sf_Cg>NDAK-^/f-g.Wf1d_^367]
RHP:47=KJXI=<JO=e2@Y.W9]/[fBXQdNT@=11Q_3)G@U-XVNYJ7(1Y)<[d>QW(&2
W12@:-O]-U7?&((J.FRF6=Y-dIdWfX,BQEbZ0@)V8HL^g_CCcdFU<gJ/?DII[34B
N^G]ZEg+6eWZ.CS7b;4;S&&JH?:\5YVMDZ&?P7+NI:8)L7SR10VAS7N#=YcGefg1
:?:dA><C]S3=G36\UNM.fMBQ;,II.^84Z#@cWR9LF[)a0Y65+GL\FD=5C3(]14He
S<Qg]>P)CV.>a10E6AI4_W=>.EN?M,.bG4fJ@5&(2^BZ7fZ1PC/P54OB;40R+(LM
&bP=F]G#U,=ga2@#CbI2[#H6/eMZ>c?3YBR>E@.@Q&CTWTC7HD<gEOKI/bd+7fH.
CF@G&e_&B30ZCUT9EL?C,-ZGf>afKPGOUP^1D81,NW941PCN&0[UZ&+B/&Za&>1[
3VY3fcQ5,#<5c)#SaF=URPQb)Bb-Qb6F\&[96MN4T8KUIRaAdSF^<\RO+ZdX__?L
&X&@EBPG-5]=BI>&9IVZD5d3aQ-bPUe:369(UCD5;@7f>G2Bb3N3AI)U>fXCRSY9
_6a#gc9[76ecKR0aL.:?gP@U+1:]bJ5_<fIR]Lf65cJ7@5((4&PZVL;_\<=&/&(]
d<aOFS5:7CWG^_<8C9fV0OTO&^UI/Z@8<X==#f\CZ<F15_C?R_ZdQ4g@8<<Q_QgO
a-cDY-4Fcc&G^P=))J\>;cPg2G2=GP3^F;H-8+a_LA]2.S)<.>J#U4),MV](R63-
0@d?VdN-;ZU,3--\N8<GcgLM-M_&HNO9#KeOB)JNX3f7GP/9,@GT(<\/3X+__Lc,
.33Fee/1YMGEXc+b3:(^b[99UgC\5G6])c<\@UDMR9.:TV1cG[&V0Q]/5[2S_KVZ
VX)1TZ@G/2S5RM5IAQ:U@A<=52^HcE5XY#F4=AD\C)?]aZ-GfdSNJ#&3gbXHN?^0
U)6ddaX/VM50N_aF.5,(2>M=:@-3I\DgZeF<@PIbBdQND)30Ea0-H>7YT_G2GAET
dU4#2@-I6\#T+5=3_0Vf<bWd]059QBb+f.-.=<B=Fd\FV9<ZR+^F^9(>N\Y4-HQ+
T]2eVOJR,[]2Kf8C-5)PH8>CH.S=(31MA#cE=+XIM(2c+;bW:\c.Z08a3F;Q=Ved
7D.@(/D0Q?FH,?SEd@&&&VH,(aM[KV@QZALfFgNd@G_RY8aNT\@c]GV@#LD<+:UI
+8M#.N._-.><T4Da<;<YRT6;eLQ@e3&RT>e+KcfaUM?a;55aDb@]fe>/WMA5QXE5
3POUBQRQ[-/H^/57??@GG/O;g(@QL28?RB1<GgFPCNT4-a_AfCM+YK#C(5L];bG:
[A<YL,gX64N@fG=.eSL-)(Cb83P7&>dPC)A79E9(G;bKB>[VOO1AD7J^ZKAYKFGG
S-4c<4)NY#]^KIKU,T>C:;W)FF31aF#a,(d,L389_B3M/Ue[eU=#Ff<@>/7VL2.2
0DfcWG/Y:G^e/Y(,)NLH7F07WJ4SX=.#P5\#R3V>]]I0@a56?@>HKVOS>:AS6?:#
X_)7K82f-)8]28)HQ&YX\S[44g34K65UaeG#\^SVF/a.SaMQ6Kg10d509Y02FOfL
\2;DF22)4Jg)^M+/)T^<F_:7O51VI^ZCS=#-&#FXGD-:LDc;&Q[,+S36=:&(eJZ2
GI,Z2gdN[^5-bD45;.eOaUeWIH0@^FYMKRc7&Z\PcDUTVE3I.WU8V@_=W:Yg9#E<
:[@a>SdQ;GV:L:HO[8dHPfB3[,))2NZ&AX\@D^.CO:8UPHf6&YRCBYQbW].+AI6,
MfR2afA6WR(=EF<2cb3PW9Re:S&#(_d1.;-;GSJG@L@;K)f9BSZ1#1:#D@7C/_XZ
7]:(EU17E6dLE]Y4EO9AUbML=]CZK-LcT20<<]1KJF7g8;UGH]PNXLQ?#G4DRd-=
_Kg;N[X_DV.a.c_QTWcFMB:a)0#<b5L=,PW[M[E?DcL9EP(E&IT_e25J<#K,Z=#C
8[OdC_SSbWRF=e86gT#V&55PG.,Q5fca13)F_#15OU.gJTNQd=-cF6QR9T[CTMF:
:H5<0W9FU<aC2X^,&EQS:4^]<)1B/G/Q_\6)]M1L6:@bSTHf\V;C.2RUY6:CEUg&
MTTI:D_b+5ZBD4K.I&Q<K:DQf?\bTX(e9/6IDX1.L;BR3eBZPgR_DYL&H=@4dL]N
C2aGS;0#246B&A^)M29WFKN2ZE?_;#6H)/9,9g]e@fONg0JCRefZT6C^6THfWU1A
7VW/c@CDc^Wc4PZf_JfS,#b-P@,dDWKGT/bAfc20P\-<1L;D\GX#]R5Of)/+7SB0
eOb^Y7c55<\(5K;52e7#+12.F_O0<4T@;;=V7J@T_+?&<7(-YKN7>5K&R?64dKdD
I@-daZ]XXQ/c<>:SS4C6-bAf7))d.R)1KOJ]8DY/cK:/D8ZYR<f,WY\Xf#;f]:G6
678THIGM)UAb/>f7(PV)HdJ5=#0aY]ce/)6866EcICM+gDKYL++J]Zg]HOd:H4CD
[\gM>(BUS&B74A<NCDE8/BH;N3@W_=4/T+;&[S86@LDafXJgI7Y&gY9aUaK;8_<3
9#^&L_^\<]<6aCGKMT@J<EC[59LaQDS-)O(E=UIV^2NVJg/P.O(M2Cg=4:UggNWF
>XKZZ97H)W\E-_+LR#M8AI]1e#<X]U=-91W0+1.@P^N;Y;])4?_#;3I-^C0fc#A/
N)AG(@;Xd2@eA)d@C)NKcBgd=K5[TGCF@#YK4g(1b9.C<_=UIG&/c&RaHL]^9PE@
QZ+G-P=KMb0cHDe+AL5)G19.,9]V[LV@WEbZRMAKD5fT,EH72-94Ud@#aV9+A=R1
D>>-O^9b0KGgK.,]X4[69]E1DM.cWedgO.&]9U=-OFDSJ,CO9Y(U@>[]M@_6#EGb
Re;@N]DQQE9F^#&&7H4<#Td3a5X2D,c0YA2S&^@:?@GTML.6+QN&BYW82#TIG>:B
8SQ-CSQI1;McMBV^LSCPaGb<27D3X)A&X_ZN8]BfI,@D0:QC:6#_@&&#]>\1?KQB
NEV2QG]SQ28/5:UgZS[.2NG81a,9G]7WHXU#eZN,9N(7F]Z9d):WCF#O:ZX<MH]0
f#ATWJX-,5J5cK9fI0f]bbe(\.aM0;&&_=YPBWE;=\YHQKI@_=68gCVfg=)(0H3b
C=6JaP>GUG<Y;LZ)-1Q]WU;.,+8[0V&F[N3G?\+CX8IZ/.cY1+A<O\[4TXaI;WDf
Q#?aFG-fR)JN+4Z4>Tf(O:\S5f]dRHYFQKKY)3\3Z.4LZ@9)W(\HZg&J\GeaI9:d
-H425b?UY0_A2Qb[9-3INHYO:W4fb8Q\HEP-VOC=G\68\/)\@.M];6)XLV@@#+gQ
THcbeE;=/I,=SZN)3.K[\C.B;:H_&H-GYFb=8eHUMd/We-2;3Q/<6Z:.,6+7<\Jf
_+[<2G70eSKJTK<I-b/;,&(_Pf8JA>::7</4XLge?f<59G;gIA#R].?P2P#VH&DH
NA/ZVN_60eD,F0[A:If(3##WGGU?Wf]R)MW:O<4\LD5JZN1P=-Z9Le@(JO\]AfU[
c(d9ac/KP/?O(#?_<EX\3b2<be]>0;DB=e8<S/e30H3?1(E)XUK528[U-]@;bdA8
4Q1B\1Be9O[R[DCQa6QQ?:LOXWDOTdEU&VXJa_9@XHc9?H=[0E7F5Pa:d7LCBOW-
L(NKF#R\#11F?Nf_KREH\fWJ-FSc]#);gTWH-D86X#P([.O?))Hc@,N=U<L;\#e;
-&C:7&&d@GR2@QN0MFg9VRB-IFOMfD5f7HSf,&,12EZTA6+g:3GL].JVYCEVZbde
ZD3WFI8OA;Q=+C#2FE.5NDXR+g)U[<[PO5OBC829Q,,G-F\P.AV5Y9&Q7-#c2UAC
)7Z00d([P_^FP#SP,0PX<Tfa;[aa2J^+\.MK;Jc=GSES>)2X(?2dY_^8c_BOZPb^
OgPSS1bKX1>G&>@g;H2(S9:HF;3:,.?C.BPEF:]FC8\E1Q)(RD[Cb,3<YSQ[=KL5
@]0F1,BX]\=1WA33+\E;84DB-X[P))[0]WbR1V30cH#Xd._N?;R9PY.U[S:T0?3&
]fJZa?fD;3]cG0(1f0g>9f1\/ST=aLS_FfG<U45#eDI0-&[IfAE>?f,WHR>\H^\E
ZF=03)L?\V61JNEg/eSc?G_7SYe?NSIWU:+9B\:+(<M0FYa<6J9=b<FBL>gFHVB1
Ib9EdBac[(1\+&f:HGaY&gX;E\GXE\S:&9BL4K]JVN88IG=b_22>1P81:\YMX<UK
C)8Ze3>(.22?#1]eQ1,2</^5bYH;BLR\^.Y<eaZ\XKI8+9b5W\IE/5Wd8.ONI2EP
7.S/_AZZ0<bVNZfI2-c37V,=]d]a2=aCL9_1N5[2WY=^QDN,c]JYfG2,@QcZ\-2W
LT1)O(UKABRQJ+P)aY&fYTWA.+LX9f2_ZJ#_:\+;;,d5ID]a(]B-WKaA2f4P8@8W
R.;[e)S-Hf7#)&]CY337=7d/D)@W(M1POUdRPT5cRV]9<3Yf4,f@.9)U9(+,58G4
<I[H/O[SDMAZQ(S7^Z27:3;&ZF7S8D-6GcUaM)7/CMDNaId4>YeO@>/N[4T#f)9I
UR(gXJ&E)F7J?<;b4>P_G0X1C)UNA+.7CPA<&F>GL^a[_+;>:800^=7S_1\\a/QY
8g)#CfLb-.MIT--\G7A7a)9FU.K9=fCG_\8P;8A1L&Bbd(5<?.W[#FaG<\L<_;DV
5Y@LZ<W.6,2/=)9KM]@:/fTDFJ^N@^P7Q=WS+4.\f/JTYG>Z3Q-),#O6\-4XCO^D
f8L\T,5T[VKdFJ^KH+T@3J-_,RDU7Za4L-((;;LP8B+13>/D>50DC3H-^U/:D=_\
Z5TIW;+C>2Z04CNA?;U0Yg^>#O03.OS7Z2>,gB^#^<ARZ+_5:>BW@THNS7faH.N6
)0UV)&XP4/^B+=&6+KIY&@+(]:dXSS<dGG^3]\\G>EeN,XAPRKT_+]@K0VbX2UEG
VfdJO9U^gc.ScUX>aBKN=c[C0=P1RC)LbV)9MMP6c3d&(K767&3a5?BZI2d^&3M6
#>99VLFODO-R\&CFSU(LAH)_N>WOT;+Y7f3M)b5/_P9B>I&.fO^Y/64g[RS,g3B?
,K0UI8YI&^5P[\RGRM<71H7+6b/5TW>K8@6XL.Mc\/Z1)E=Wc:Y7#5XJKZ\Tabe3
T)U,\JISTPG54_[/-d;Q@1&S;A/T>QD3M<RF6U@RBTNTROAg+;ODYABga_2c)I8J
810C_=c<7EMDD=L39K:7-7FZO1<+)\dIB.P3aJ36GB/LBL\f<QW9;=;GY76Vc\)1
ES_&?K&RAF?FXb9BJ\6OX5>:.Je#cH,L?VF0,<aB0f8R?GKJVN#5.A10[2f5#:P(
T#[,8B^=]0QVg(4Y4a6I9.XUgd7CR&I>5^L6&<Y,W[09J8[,.RGbK)J\1c8NCZG+
VMCX(706M0>&aV[[.f5<M_#84,A2-a,fGB4M_0K[f(c9:79)aZ98acAF]_186[W-
ME_V?1:9RN)bMI02EcNQ57)5TKR?9\&gC3X]?=&4.]f;?4M.?I7@&;QR9BP:P]bG
<Y3X<0_E>_dcg1/^I_Y1J;Y-XDg5/4[Ue:?#V[.a0CVC4L8A4;6fC(QORC<fe]#P
<,?UacL;QMB,A&/:BV0Wb[9=>PT0NZ4[G_AZ.BBSN?ebg_e61VeNB+2V4^cfIK-V
Z/f?L6?;)NdcdJMaeJ?_]31R)cPP/I4;966FeLJ21bc\:7c-eCT3TVF3a7Uf\Z;4
d&c)VJ?QU:K_A1#&I8X6E#P07D#POY54GGb_FG:;2:D)Oc0eF8<27W^Z+LO0->XX
f\(=?d-[+OEM6-c7)Z.&.55KNcNL;=+XbT-G12,JIFQ_7I[f.EHRPUKNVA2Z0LdY
C+SHK]>1LCDZNZ[aFM;M05;L<YC<E]-#cM9<.;6MYbS5&T#E_+&E-_Z67EL1-)JH
9Y8)Y<:EY(]SOK5S?;BF^(>QF;01\712^Z60=YNOc<S@.F\F3_g83W57QFL;FP/g
;Z47\S9PW6:aaA+]9<R5-bcNUYHGP//JDEP(GAJEN9Yc4;7Yc>H.b^<W<R1f;XZJ
LKR4TK;((^Vc<.R:d+SQ#QQ@\+4+H864?G-0IV+N;?8]^SG?@;\;.N9=^&8dYF9[
ga3fSJfWR2IbM6;39\#9>@8QDPaMFGZAV)&J?_\\MH&d1eWfb)U+A@9(0/ZOPb55
T35=V0P#Z3D/=RT1+GZf^RO4T<GX49P,@DXV^Z8PU(()0E9)?7I_?N.-gB8-fbRX
BF&c<_^gg#V,b>V30;7ODB1HWH-)I[eH;Q_<e;QQX[B?ZC(/&?Qf4,N20?SZIIZ:
26P<M>+;MY:+Q?(CYRb9J8(I?eT,UMTZ+9=+Je8HKN1=\HM@2L8I6:F#G[(-/4[9
Q/EY>D;7]X1]D0Z90I3@_SON/^MTK&-;Eg+8HdSfQY8_GdE^agZKKRP5L:T&IIOV
)HIc9Rc,.K4bYBdd_/a5FGaN.fV[9Y=]=U=1U0(V]NCZ[@DTHD=UNUJP+XX]+UH7
_8P.A/,=:;7D=LHQLF<H:@C0BR]aVXFN1T7->P)?ED]EdZ;:W;8&DPKBE//.)5La
f\H9]@.X+5G1_+OO]85V^VN,c+D8/XN(8T?[>MEdT0_Y^/^H.&g.RY9:-#@V;cCU
/O)M6^RVQXRG+5[0E5-a;:ee-C//5GSGVZ\b@Z4DZGfD31UWc8\GOHW]#DWWfRC@
Oa8ZHKBX3?<P7@0U\R+g0ZSZfL5CGH/#8:4FMbX[,MJ^0b2R0d&A4G^P316M[eBJ
a^LCE[.FfL^,@4GK?H[R-1dN]4RRfGS&4cX^B?Kb0A,D];#[Q()/O?+GV&H7A9B0
>]KB_b&TX22E57(AJ@F;a:cedWPfUG#Q6LCEQ?J]1#RU1O1Af-A:AZKba\H.FD[_
S@92>L]&^;@;PU,?,Z055FU:I4M@=WRT]\5&K17dV4ae&eDaY2cUeaVOIOE3;@K9
98S^@/:8>O]b6Da&O7\KF/VIPX>V6Ff#7IA,DJ)<)6_[5KY3G-?#Mf/Xc[6Q@50<
1ZR\?adWP]?_]=9RUY\39E.]_5BXN7HSH3_]P(<CO9V;F8eK:FV_-CK\UVY@75VP
E(PR?QVI;7ZFb/D&P:FHH#?1,@f6I>G/PbJ1KU2\WFF@C;E<1F\cM2aId\F/T<Sc
CS<IN)E[0[(&QbR:UEN&:Me,Q)95@R,b;D&T.#70:_XPS,9eCb-5-g=Z-@V\\YE0
>5g@DTF9IcHOfD<N;#PT<^KPUUVLa[MJ;Da#LT9CN+Ne0DgFSU(\KQQHH@GW:EK&
IA^(SDTaN+V-HPX4J(8]0@0.g+@K#;#HSAdV7^>;&0059@SUY=>H;0S99>;^5#Tb
)D=IG:FQX\O3-5>\72UK))K@[U54B6^WU0#/E]VA6^#OW:WJSdgW#VISX[&6IX37
0TCC(LN+<;?_71VE1N3(MM)eW0aL,&R6XIX48FI@;/)d\V#R7O(2+V#XM+<g,gX<
McI4IW.\?]F55O^N.=)A):YW3E<Dcaf1gf+]:ELgWLT-D]8e@VK&RQI1GHOKWC@P
8QHF;a[;-OT:/>.&>R]ZSbe0/8?E.8g29b[]e8S-@<#JA&=dcAE^fY=]G3;>P>GD
?EQ2_ONbYG39/Ta#RZZ2.EZ/PM(GgeA5R1g6eM,5]HNfRT_97@eRH8_?K<g9X9f#
5ce0;P4JD]H@#be]8(,4-.?3KK:+DA(>R5^dBf+>+NdT@@824W)?B,.^CZZS(gf.
X(Z7KIZ^gfZbJYZ-./(c&c><27\J2+b2^P++J0;SG_UE\MTMbJGFXQAR7E7^J4f-
g8XND^_fVA\#@)Bdf7E&H]YAM\F]38aHJE-WS>5X0FWH=]:@?FaTF?,<Rf@=I[b:
ZA7g&KYC#,985ObR,&(cbg5^S5(C][eT#R5IQ-P#M7[:A9]=&>0&EO&H>e^=gc_X
KEX,?2&X^f1-+g=:)/PFPM]GEd&&QJ/&&4gdA(EdMRb]T_=83(eLA?ZQLd?Z]X-.
/O\):(f?PDW^EE5Zg9]6f2K=:CO[OfD>2LT/2g)63PE90dH&E0Q514Ue#8Z11da.
cOOMMd9RU+KL6QEF3d<0@U6MTYD-:[[6H^5:F-7N/c(a0E_AD?BSB8Z(c+)M_<3P
U[D46b^3#_2P?76X^OQDb>02P]7:>Z4e=G=HAZbL;RC(^218KdgD>5(@ae=:_0f/
b-e<@Pc7=/@#&UJW.##B[&-Z;EfK^&WF/MH/=915GWad<=AM]bA/ZSOV/[bXCE.K
()Y-f0Y4Q88/F@V&(?dS&gT2L[18g=F()3-BT70Z>>H-J?()V8,Z-0D5-]A@A5_S
BOedYMfEb5a<B8e?:G2FH0GMU)HO5e=Z]FbaDfLJ?BLVb-dOQHFUNB+,M<6X<Be/
U;F[RLA9>Sc9Z7F+F9IPTeQHB>gCS9@D1<fMIJ?7+)0/+gZC/d7R:/=#4P^&5PbN
H#JUb=)[>T#I79I#CORd6@c,gfa0F^.\(g36G^d5W6@1Z7.R=-LD41)H=ef?,=61
PBc7\6D9dP0V09-K]/KF[FZ_Zg=UTEE[AZ8db[AIHTGUB<62[?>0HFCY9F1(9YbS
AY9E=gcRg-J@^,GODZA.5g[KG.BS;#UV5fIW8>/H(-<S.F@,=MD#g)4;?>.-SM86
3VI-R0VgZ:1RPM1[f,Ge5<Y,/&I1JUZ[U6<O7<M#;WBAL-feAV+6bU?L#;=MDFD_
-+M2G;.?@#@X\[5XaYdXcf.WD[K;5Ie,-;M1dWYG2LDKR6-ICbeJ\0JK#6_>([2F
+<O3WaQL[)SLUadWb_#,OU.VA;K:>^3e0_93Q)^<#efJGJ1]f(/LCT3[NJZ?>S2.
WU08>FC?gLQ;BUIQON5N:d5##WH)2-,<FD-C5[Hc(E+37XLN(9&;C&^,B(B#0d)L
B56SG7-\6YH23--V2@dg&H3Ea<:Yda,MX6XE<3FZ7L7Jg>eLI26R-;)#/PG#;XS]
dO,;_K)aa_]a3@V#CI879BJEe6E\71D^E?J]H7BP=#f]D&\IML]AB(:9^gTH4g1f
a50N;P&A7aQf(^1:-WA5ZEA(eF(\-9Hf>22P>K1+,6Hb#NCZG;(Lf:?:@20)/GEc
JQ75c8;\+,g;#.2Y0f0g&0cA&]@JPg6Z>S&GZeg;<8X>c]/5Q^?-]L+e\b_a/9;:
[^8=gB]f1<A_.?@cBRG#;eR.cFK>^<C@/I];<GJ9ee)H(daVOZAMLNL90D55c>WG
YM^YQPV#SV9JO^BVR9UY053J^De\aDd)>4J7ZQf+C_Hg48QO33cEe?f+M.Z;63Ke
TX)b/C56e\RI\.1T-Y.a(X14L#gI-W5AO.\)TO.#d3(SPZZDM^ZML;7SeDNW?NbN
R1g-ZccTHL]7bbTg4OU9UO44DXG+)X\FBc-HQ(OT7<FaUGTM@65[VN]F>2@HYDa9
L&c?Ag,\_a7-50Se=LWEU,N_2F7<#<]-6X@3QGH?L?+DW_2CT8bDQ,@D1JJ<=8/M
4GKQ6JXgE2F9bE0b&d#R&;7QRC-E5&:/GSOR7K^?T1Ce8J1cAQfFHE17Tfe@C03B
d3ARL<d_L&Q#JPY6Z.?VI;.+#gdY2SV<)5EcUVTZXaC2L(eTRU9A),XC(bRY5XH:
bVbU7Jf-Z&cC>^a/O.fdgP,cZ7.>G92Y=3SE#H3YcDO.[Y3=6I/Gb]&=4QVQHIDa
L4Z;F7^S(>dJ0gJ[<Q9g]_<&>Jec7Ob_S<=01>:bS9(<BAb\OGOg;__4[1SP6O36
7NFC+6ZJ5Z=3F>-(&8R?Cf&>S6WUe;?HI.7>_XbdbbgX(04G5S^KCWDZ#f)6Ud25
@J\a8<J#a/c=bUUHR1O2NV^^A>RSRU_F_g.N<JXf#b]F+M0G=BQU^O2IM]KYHag.
^F[EKOZ#W]>-=^<D2eD510#.J[XFC^-+a-(<D2Z<:RHF=[N:Fb:/N,SN3^\NQ0f1
\)ZF;GW]eX5Y6ICNM6M,Le2V8d@O7-M,-&ILRDf)<5EVaW8HJJ(I)\]UJbd66Y=#
X(]K[BRH>9:g-,Vb9=d8J;Q2YQO)GFURCYa-._=eKMXDV.a80:?#XDW>KN]M?YOU
JEe#N5?]:cRXZXf;[H-e?F5@:Y3H&cK0UHcBR/g8d<?/;+GIE68T1@bdHO(O8WQ1
(A9JBYO82LSE&1#5>Z1cBf(I3P=E:IJJ\,.3QYE@A_fQJFG1(RCH0,L2#:c\2_C?
UMMKMFZ6[^dWN\^+T6S#0F,dMF6]dN2N08SH8HE:g/H(OW(dHJ2[^GB)/fdCW2U7
:ac=EVMW5;>0.dAQgAS50aJ:Ca,#N00MfX#ZaE&GHf4>2^L.QV^[>G:##GO0g=)c
X\CDQZgSH;9O>Ee?[=9Mc[TDc9Q>@d_B8AcE/Ld96\-LIM4S++/#V,TM&J]RaYe?
X7;SbGU_Q5,9N0BeI,#+XI/;:]e-GJC=La260^d.,X>>eA-6aL6bfFbZ@PgL<IJW
d6Le[<S;W7DS<IOU52c)+RgEQaS9TBDVF,<KBV7&_EBLL#37_:R0Q,cP(-#@>gA)
[&K0/d[KEAE5.cW]L=&G^+^<RA@.>[._;Wg=9+M-gDJ:e[.4N@[>&^]HXb]g-\)O
eNS6OK.@c(bYWD2Gd.gJW7cL2Eb4Q[VL-6#E>1>ZTO-=M0[H)UM-,61S/bHGJD\N
5FL&L/8ee+1^5P;KH#Z1.-CB5eN=358\X/N&ATM=)T9&/NS3+EdI]L1EHQ8<_/;T
a8.LAIF4C+/>egN/[L[R4b](F<7/7G[44Z8W9]F1bF)NK@c70bDeR;3[EUG9I;/)
I_b7,Y8J=?:&\W@WG]7c]Q)^E,&/1EMP-La89-[:2VFR;G84T1ZP:X9Q)NVM>#OO
-=AK+&[U;c#Yc_E=.#./Z5VOM@HS@b+P_VI?M9R/B^3f((O19^U<_;-cDT,I<L<.
a),ZQ1g?3MP0=T05)e3Qg3M@U103#7?0bT:DO@\@0^)3,F(gTB9)<M^&?3<2X67(
NS1[7H+@+/CRD6S9gOfSDX5^1V?V1O]b9/.N3PSO07g3V_CcdGW]g4-2:5N&AYC#
=c;>d@)[19A@/g2[NF97HUG^=gVG5Pg0Kd-?[(&-4RNQW)V_ZO+VUc2_4^J1e4;b
f(H87)G^V9APAg;N2MAbFTCK>>>9Md@8Z&8PPT/e=_dUN8&36C^Lf2D0<Q:<2If6
Bc6f>+UE4^aP8]E@#9G2gA/dF-71TEgP;EW7IME[MTE-#GG:C,CIL7a)M9AUI/_&
]A7NN_]1(7I<IE;;M;GfPQ]DPKD+:#Me:[9\aKN,RZH[MD:GR)=.>D.#REV;2]A1
H+I[]TJ@MA#Ld\H#T?/V](Qf^J^/4/Le9g[-/O\XY2>?VdaYN4Uf9Ee]=NE7_5g<
e:B>E386NBd3TE;&#4S(@.2I=#@V\Ie4STC8<E7H(X^]<<^3HEDC65GdEM]=@ea?
?0+f8.@7^Y>@^2N+VQM/N0B<b/4UZEBA/70ZAa)YUR)e57UO6a&g\/Z,P@2Q@f0X
WAK,;-M[5;/-4LFC3Q-8b/Ma>0MYSX,GY.+>RIUC<VI^8GQ<_Z2\EY89d2@F@&E6
(4eH6B6\BEfRCS9bW/WTeT<[ff)NC1-M5\?R58NfXK^.4M2K3LVI_fc6Ld4]C^<1
>?M+;8(#S9=?cSNK6\;G;X1Gda.\&,4ND_&S4F2BAKOD9CZSB_cdJ_82EK/;5#72
W#3SE1]IAeVd+]Y61aDCBOd_S?J#)CLLfcd?BXSPI>UMGHD4@/>P1NBYe/#,aT+2
JU#93CG0SND2U^82E^VIeG]1>-,B9/BeOME8D;#Vf-.Y:FOb8F;L;?S&O[f1(&Q8
E2=[S_4E3J35_(d26aU@&>J>SRZF&DDTaA1:6-[I6:])OCY5>?[]<E-;EUE5Qf]L
==K0;Z5K?HX]K4PcJ+CM1.SPZ8KKLO--X\^N.fI@:@F@d@[^=eLJCKd?>3W)>J_)
(L?bbL78>.GAEf+6G+,:[Zb-e\-3:NHF4=1][NHU6=g4R_d2:\9&](,H#C/M..0.
D>RgHPP>Xa)ST;_R@Ef(GH^g,G3bR4>(fR=FUAfOJG>U/W&g4&##.V5=E:XQ:^=Q
S;AT,GH09O24LSN15YG=F6UOKf0?[PVf-H:ZN=Q6Q[NAC+5YBF07>B:C[6E4Q?Z?
<MY]=EYJ7e0S8X4DVGND/SNKFB_2E_K<1//56YNIV[fd0Fa1W]II81Jc[TR3O@[B
NG@T&WBb10=f7bB;<ba3ABgd=#FH^\E?V?f1Eec:SBcM30.6TO5<4([EX#94/8_1
R1.7Z\FULg&;TVYOKQ^@\a+G/SPCEcF>\(YbN2[9MPOf[dHd1VQP0D+I&+6[(QG]
@XH+,6eAfDbF0AHaV(dEZCZC(87.=H7N6I_g\U82&WFS#g84HG7A,AWd,H]aALGd
23?+<9N1LNG4Igf8^@/@O(Qbc&#CR/>C-)@b870XgJVd;YY<5IC@)YD,3La@dY9&
U+4:.WeNOZ,?L#.<D^V+U+</IFCcX)d]:fP0F[Y1Ne(B;PMT#A4>?^+,fWY[V_;Q
I(Ub/OFN?/(J?730#cBTB(GgGB+<T^9Y?;)N3(TUGgW0dXJ5\7&X.MC4);N_fD,6
5B8#T?eN>C;YeI9/\a.6/7AOCF<Dg#TPe/P1eD]e<M0L;b\cFF1Cf^1<Pe##4VF_
G-\?:.;PG?@N<@TfENa(38;ObL5>&(]2=C@,913+#KSAK9&.]<3T4Q?IF+_=S;H\
<J<f9SIa&VIf_.L-^]U([-.[E/:<_:@4E=6H^\egM&g3R;VYN\;NJ4.Kf89ANP]#
5)W(4EUZYN;a?9)LEBDE<]_c#FJf7aa_XUJWS98(g+#cba1MAeLB,(TReagF^WYT
5IUBLO&:BH93//&YC\a,9#Y8;+J+Z5EJc.F,T&C;QREKQ5:c&eQ?7R9J>d]Z4UIU
Rd)00UI;9,)L1P2.;>F(5&H6+R5:&f<bI7/[EGGLDZ&B25=:G<?XX0#]VRg#RCLN
2&[J<ZXg:e&O/,a0XW-d,)NAN[JDga=FYS[@^^bEF4SO[2K8J&W_?J5NFLLaI1,c
La4=ZIb<GQZ<;LCMVU#T&]ZYbGMc/4I-TL4/F[-RX.-c)Y[BC,09WaJBERNRT)GV
(CBbTQ<cK??EP+;#QGR0+AgILa7MO(,>AE?e=9Q4<G(9#IPaIJW,KaZAKYM[<]45
bO6)SW<)cGL5D3@Q?f3;R\RSBHF7F2S1,R5(J6c],]8=\H=EHP3Z7P]5EY-?.,gW
I[Q38A1-HDPPA5S:T8^>CLSM_:I-CcIUG@#0K,6(WPbbMRT,8c=U9N?UGA.U@NNS
2];ERZ=3AV[4V[ZFY3<B=,J\G,4RV/0=/K[#4>V1P,#e#&=[d&-BBf#;]BX#=G;.
Z1S>NWPbg_1aY#I1Wag^\+GIL,Qg;QNK2Ie^:d5[1GLOX+(+:>RWG-VJ,D6a@Kec
L3I&VegER>3FHRB:WH>b3B_G=D@^4OMFF7BeH&B?D>1^WUY?Z-6Q^CA:_,L[UHRa
ZRWD\d1DW&.][=6\K5MND[K8<&T0Y.Ug2V6NFQQV/\YW?ZT3:5C;?I\b\ZAB&=L)
22]gT5FS+BOQ4^2GEc63Y>,K+cJ>5B]g<X5cWJRC-;M)Md;R3\]D5^_]F.&W0P9U
(&acT-e9^8VNeHXD)ID)QBT=/PV9,&BNE\/:&S=?QDLBUJZS4#CfVZEX+7/N6AI]
4gKCRe6-@E6S)>WK8>X#8\T&Nd/bN1J^7@4)N?S&BC\EfZ@&H_-ceE7,D6QQO)H^
>B]\Z;eF(e37_][#6@A?c?,T3L)]ZTLbY-QND.86&gd90RUgGS(W:R)JY@ZBHG0Y
H#08H[g>N48Ldb;bI4.&dg\9:+^M0_ZX9Kf.+2W:97(2U2ZG-W7MIL9Z@1=9cUJ@
[I8eO#32<5Q,Cf2RQF9KJ)Y;8aVY0cHTW68]c7;JUfPFeb/e<.K[URfB2EPN@b52
YE6M^6S4WR@,J^E>-\P)+IB839KOb<Y_S;([@5S[DN@^&Z[/cW]&b;,)AHQ+d)a-
a4+PW_G-&P#CWJ5IFPG<.87MMGC-P4c0Z0FgS@MZ9\C&I=;@)?+e.8#+W1SW<f6V
NUOTc.8T>1VU^O8:d]ZUM=.)dPAA<gQ9WcOgYQAb3HKES0Af(/CccRb/5gHKWY[-
d#VaZXbaFcESb&eg&>6M93\b50&0e&EB:_f0T_?;T>:AI[]I@ZFeHg9,AURE1QY3
+XD1:80_;BM&.&0L;daaD\.[SQ_UaZ4S;E4XHN>>].4,/?+#FTa?K1H:KFO[gQEE
(TU1_2=d8cHT@W?fdVB&Y6&XS8P+dR3.M/LI9a[I=TWA@YMGF;#<8b3U-J]O=UBQ
\A2H/TXJ_-FVVdB#+XH\8?B1]^UaR#a)f<4B3GV)@(KAcN.UA-LQ,&43Y6V7\0:)
be=Hg09<QU]U>eB[X87PgB&GYTZRB@\6+8<TUC2^O&V^E@AO9(?d2&G@1AQWM\EE
P:#:/c6d0@1TG>^UY42Y_<6?E=5fH:P^;+W/9?U]BP+Y\MVD6G&,V,/N2QF8:@]g
Z^K4@0_A<)N2S#/I(7Z/=,/EQ>-T)5/T^05^NgT#-D0KKG9+3GSaF^dEW,12SP?A
UOa3e_fUO<=gS4SG@8bD]=\Y/fea[[)GKMH#]\b)X<f)/?KZ@EQE95V8)L[4>[H/
Vd0Y?J]Je-\WQ0J1)L4:]),gSgbATd@gB;QcOe0F9d1KTFM<0WWBK=(LTC_dG?/\
LZ.4(?+K)7g;+1e^T,+,^4RW30>#L]I[1N-87&MYR4@UBX\D2D)TQ?YE?XA4A<Y@
+gQ_WXdXF2V&.AT_>3.&2f^OJIgG]BF1(D:SMGSO;7H.=?1:]OTL_F^FUW0I9&1A
#<G8Ng=[#dBM^VaGb7f5QODdPd4):BA]G-g>XP6,_.+3F70G@G/697(5EUgZKBK)
&>+9_Z8A4,_H]I1WS(@O9/PbC<b2RBN6ISKD,YL,bR;FHB+V9TEO6GO[SDZ:Vc0\
L4LGR3VYRb7f#E1ZJ>e=9/9[M-#KNL9>3^7adD2:)FbC?BCBL57PIb<\W/ULD73X
e1bL2@CfY=3_gNXGGHC:Q0P=C6UY0P:1f[[GKbU:8Z=04P0ID_(=#;<WCW/b5KQ;
?GL]Fa([bW6L.B2\Rg]F+c/.A1))XMN139b;;2fV&>WMC&?657FK(YAI?_5NJN=>
(/D5b<Sbg(cED7Y6XdfP9F8.L6QZFOWUYbX)5935f4C-S1,[12;MFM4>,Nb8X^B\
eV8[gRA_LH9gA=]N+X8-&K7^eI#4H.:f:S.#Db;FVd@W;C@\PXgGVW#J@^@1-/b4
MIC?SS4C3bWL_Ab4EgTM;C[:P_cF]HCO_KT):6UU/gBQMSF+\WQ]7,9KLE:,Za<K
d?.B/1S\/T<T[Z1Ea6^;Z;_[b00UfIG#2/GD2^^3V+\b2M3SYMV#(7_eb[TTaGU/
YT1Ne8+R<VL&[@XX4b,I7N;WdPA2>X6^fcZ+7;-d9\WINAMNe:AE[(?G)^59CIC=
)NO^C10W7.3&D3(7.N<I>(MA&.:4X),676;_GUD5N@NB9^GZ9&9K64IH3PG&5/,?
ga6\b-SgTA->+B\OQTK0e:)A;D:1[g&.>[)_ff9CSb1]+J<7c?GI,/Z\/:(YbN[C
B&0LP/13:_-E=[KbTab#SZG<TC[TCd<NF89)M0Ue4/7:2P?_CI](-dD2@-14])X7
H4\O/WJB?S>J0CF:KB[-),U1EM9BJ\+:AF4_91HYC2f^_HK/IN8=E2G:\(,gYVS(
/:;L\Y9T5+2b:Pd[aZVTQEJ.gKJ>;;8M8eb0L<0;=UW0dYA<FIc5Z>IIB9=8SE,H
N.eJ8XeDBfe/3^<J#D.P(,-\RQKCUc-SE6@Ye(AM7KM<JSVEI5LVGcQ&DUA54f17
NLBTO\-;@U^3S]:b]4R9?:]3P^0f)_+>Xd@]]bQ0(&VH^)Y]Gb&_9JVR@ZOE9]WW
cGL1(-V1JFbN0.AX6Xb\47d)JFS.Q=Y#@QK)D[[]Wg(?C0/I1C#^RDQ##cgDcfX^
-aFgAP-_?/6JAELC<E8V/.Y\<WF<M2_@6gF-N]D<AHDW.&7JAI=#2+YSS@)F15a4
S:FI89T9WAU#ND;Q/?DM+=NPB5eZda#:/^d\_@MAN^8R.VO]gR7;Hc7X8,ZQ)21D
IadK9],JRJR#CZ_/3WG;U]B+)CYFN>H:(E:FIAQ12C8Y<TI8BZBKC.UYXZ5L\a+V
@:V0g)1^CJ.4-5-E8f\(EQAcGaSJ0&A(/F0<NG#ET?-He]]ecUJU9\79XZ<H(E2[
.+315&SL_(gH/X5+=]FAFM4Pb)Y\:.D>cJ#E#ZG4F:)dJ>61^^KS<;YLJ(P5E)eB
/OCKA>KEJ]FLM,PHGAOE4MbEcJ(O#gO_8,dC9&S/5b#L&_eK@89/F6BAaN8SW_96
_aKD4]6?<@EV/JUbE+VX<G40NX93dFe@)e=^F.?3=-#:dTH,.Y6HX3:,0Z&RT+@X
/&D(QXIE05[a37.K_6#ZL5?2Cc,bC<(6+I5QX9U&3_\S\+dJM\IW5][673^e##(F
S2R9@;G6:SN\b.5J#GK;K>aY(-gdQ/?XO:(DUd\P-KS1<I9W(JUQ-5>7+<Z;FK_1
Pb1NM#@/L-cR:\0J:&2gR):L##S4]3fF4KL_UYMcVF\JBL]D\4dfdC-@]2KCND,e
@UT6^9C18II2g81;CS&@Re8NK85^a(dU-eNTD#H;]a=-0F]<3FHf-Db3G\PER.O9
bBWT5HeFS>2G:;eI4#>4;;(6gI8JOe,)]Y1YA1)g&;9f+cf0Aa]]&9N_>7gSUY0I
4&]N.JW,I8T>_6O=X2Ud476gB8?<Pa7(TSO6S.1QHDH_863K??RAaMRC-[KBLPNP
L/bX30ZFLZV8&/Q@DcW&8X@5<DG:FCKHXg7dZ5(30HA?(2Pc#<fN3&)1^a:&e>@E
fD:gR6a_e;4\7T6I_gS=Q2L/G-Fa)#-P>_#K6FC+3[^aZ).#;?_V\?_F()KD[c,P
2dHW)>CILEPISE&#b@1.C#)84TBH1OXCN@EW28/G0_TUWYHHg?U)SEUM.e.[WCMB
[L@9)J-LCSTeVDK>,+Le6^\4a#GZcXe4.d[fYOV(e^SdIJ?b[?[<9Gf8\V3L5EYQ
)&]:JJ4c&@O=QY1[9[O,T[LZ[d_A3ZD7=?5c3<K6&]KT1XR#^;J;E,Dd2JHVbgDL
2<EH\&dXD/:X#Hg+fcMg1E_D4\]>9A:PS?X9FD#aF-YO(2ALJ-.LQ-eZ0VLBFJf<
3\LOUW^4)-VK@O13Cc5RC)dI-:@1EVE3C8QSVB424)@]L7,D+;^=KOJGDN3HCSBQ
:9.OI#e:SP6^]<a_>C<_J32a+;A&a]PSJ>(S^)UZU?6U3>=(U]UJY1]-?-R9+^U&
A640[0).@fZB).1?_6W\gDPA\d5XK?W85.\:2_g1K7NP03(UVV6g,/RfP4Pc,455
V56aQd.<\Ge>daXCa+9_]+IDH)EH,eKFb.;X3+GX/>B=?FT2#\UA4Z3VIX#eb#B?
eYW@AL0)T[JJP/LBR)M&IXDa-eRfY0_#3+Y[V4?TY->e[RHXDL[^JLH-0H1U6LQf
bPQE65\>bBCUTFd+<QN4]aa>1)G]W4N#^H\3P<_:LVJ6gcQJ:2+dUE30a[ba1L+L
Y?&Z<FOUFR,X0<K#YM5GK]WF\S8/DEb\3=FcG7c/+=1VF+Q:DY\+fZ<#4T.e)I41
OPeMMM8/&M9cCDOT@8dUYBWQ;UK?G+3>dNFM;\[F[O;4^OMPPES(-2_X2+(W#OEP
SG1I]bM>)@X@;_+dF73e^].I=)e.CDIG5Y3C_e.0^Y@_F/J3fY_:gC<Z\gX)FH:P
N<QBG\G,&O3XLX;Yf9ROg]A?L1I3I_>W00g#<W/HXX,C.IBM[S@DN8]P:7-2E&<1
33RGEM;+IQWU]gPaLS9MJ<\6KDUO41:Q^0+@Qc(6:OPReH#\7f;(TWPed8CS_dX>
]gJNfE:T..?V]g0_fBdfe#\=;U-97)?S?/^3^.V9F?cEd8gY=JIK8Vb^<JXA2A]2
T/72E]eHZYGVF/HPd,V?)F#SfH9T7/(Q??gN<g[Q7D\dV;f[_RL2HI,P_LdeATX7
K&#EH7W-C]\BCL2\>:GJMPC^+R/_&SX:4/D_EW56WQQZIGQJZ>9]AfQ5CSZ4<C.Q
HTK1\V#TMT11<2N7B^C4?&3cU\Y+c[N]IEDFR?]1(8/;0#+E]I1Y,-FD-[?,aD.M
;Lc\WHPg-(+EcDT5HY,=)e&^[4(VbC?[@Q4<UQN4e7A+E9RDX)[2)QGgg?e8OC4;
DEBcFN+SFQ]9YJ5B;A<gf/E8CgdA7HQB8@-]QQ:76/CL]CMLI&e<E^SB[DT\>R&3
4E]c44J5L]=/,+R;K+<WG8V>3K0WN&-63/10g0>QTH4@;#W:A<K&N:C_0+0HC82;
E>cJ&d/7QE#B8B5C+]T\bf)aE8Y4VcP=>dFXeHdKS3YGHL?G&@?XZD?U^3/<bT)c
>HeR24(91#3b]P-Ic6X0<;+=;,gaSFQFbRcZfH.5@6ecFONXW;,KJFgEWeO3][aX
/./UP2@8,P?Y:SFFZ=4ERIFBB/IL&f_/<=dOIH82K;Wba.H/FE@beMN__=P2),.U
JVB_=B<?-@Xc<_V5cG)&[3K,FD:L\A_K,JeVYZ/DfaL:NN,25CMM+)DP=149c?&g
.\-PC5:a4QaAW]>@f[Ee1D^dgC]M0_RT[Z=#C8QV.afH@b5\V25,URN2.-_QW,03
UIJ6gI@.(bKYb;OAJ]UGf-QZafSVAfWE\^gPT6ZgN\BGP<@BFZ+;OIB\e\A3EGdE
68V0;(2,)-82U0I;AADMAUU&@I7H^.ME3OL/_28.>\Z36KF>F_B20I4PL1d@SLHK
ISc+J8<OeO#8IF=-gCLOFV^H+T=F2BgAMU71CFYA5XF4&/W/DRL(#51-K3-;K@BN
C,61]_Sg7^ZQ>(Yd&9@AfKMd<1-(=G29:/+(]U#NN\28&g(K&N0U=IC6(/9>bYF2
042eRETAS:3[AL#NO3:TWL#X-4=1SAL(>6Rf)OZf9IQYS3ISC^F=0YROCLD(XEb2
>UM&[56U]_RVM9g)OQH&b7.MC&O+=X2:JU)S2b5WOZ/=1gIbb_>;3<&\4WFVYG[V
&V4#b1eH6=KB00aO:XUVI\6d_U^&3CS?N),c+@9BQ@8CVD25^c<&XW5:fe_RY?dP
+N)F[#4.[;Xag\2GOXc1GE+OYXZ<R,W30EEd9e9VI9-?4_?WM]4&/V+]L==8-)H^
GYJV>,16>5g)(D^8SY#?5J:6_5?R3(LEF4:SdGE,<-gF997B;f29@7]9&R7;>46F
KEB_Z<GD079U(C5-G2,MgS>CVKS/Zf>2D2W\GgWcRJDEUJZ2[R>4V264N5>5>K7,
(,KO]27\&8#>Z@C20IZ94Q>&21c(a@d&b6I-+SKK<NgONC.BbZI:Z/GdT9-F;f=S
V>Sbe(WL2=\?Q1K=R-1APPV_PE@G2b91S6^c9Y)E36A-bF[Z^,]#@G0cbFa(c=S3
[#/NVa[5cR7)^f^ETg\ZV\ES#E7&7\:O4L>fV_V-:]1<^MUJI4L>8/Z6\bP@=W[&
eBWGWOZf[WSefQI.W(87;;=[&PR;H5HUU.I?<HaU,_^P9;T+TB>f,d&-49Pf0P.H
f_d]R\9;O;>F>5Q:GPb:_9ac8e0g_=P0YU6KGLRIWgA46ZM<.+0B:M^Tc)U(e+Oc
;Q98S,>LA@cKXFJ6g@@F098320VB-g?_JFL0Kf-dDXR=ge3-I][aZI)S)c#c:g);
WU\P@)NacJBSdGd^&&D]IH>SD^->f3^7@Paa7CVcOI8EdeN0c5A>=S.]3V6#.G&E
\(X&J;-F484NI,W;<H/a6VC@g[^RV0X&+OF\RG9Z^>RCI@)-Qf&Hg15\[Q+G(DgU
PM^8RZK)J9^aTg=0>GJ:\E_/^]UGSRd>PU7.F)NI1Y.EG7U[Gg&a=@I1Nd\(eR)<
N)Q+?2:F)DW/3]<E^eJf<6be4NCTZT[AOQM[T_^N&:04H\<bM9b5V1:T8E]QdC9X
g>U+c6QNGDKQ];I_D;OF=6AAZ6=#_Wg5V10NF:#/4c\[19BHA-AaM2@fgeQI,,MB
f5b)/LLY]&Bf>-SO(98&6>[-gI5bQ#Z@]FS#2HQLMcNO[SV2AgYHN&M-1;@Wf3T=
c/#9R?9<^83A2]I]_XY\cdPK^/2FDKTMe3>0\FgbPECY/HKgVZ8&.WJ=S+&OI.V0
JYcG6g\Bed^a)5U=QF75e>-4;]>9.L6d2@M]<ZCN9X@_;0>_KcKHU<TcUXCPJTHG
&MJO1^8=?8(4cJ<f2C_+):GQVB,gZS/9YYCfFO^fQ)ZERG)#b(;UgB=BaWB(B_c=
:OUXGCUS4;#6=0F&;QCC_VSQ&=S1)7+5D#KdH_69O;?e\OO=c[eI#dV\[W/>fgCE
gc&5I[6._Y^4H2KfM\BfJ^?Y_85<NB;8;;KG[D?S0V&Y59#,3B&Q0-,CYR&DK,RN
WLA2&.NHbT_-+c@QUI]aI^90+>HYE_K@DX?,.C2,D#/RBaS5:X[+&R:N^Y2W0HFA
L8g#(#EZ@,:+[MQ(VG:WN6Ge2P)&1G\C&7Jb-g.MCH/TNR[QRacdT_bT/K,0RY=K
2_DgY]=HceMUZ@X)JD;g]VK]PD7c^[=01ZJZ4SE&L#?[-5^3X6Je,<bRYMc#)aS[
3I/E5PY;5SF0B0-SIBfT_AH-;DOQM],96N+8E\YGQ=^GRbI\eST7=&74JHN)fY3&
Ff=0O??Zd@,cT3d=K8T:0G[WUXf.Y:f,701+;9PD1C?DXFdXRb1>M5Q:)D.0(#f2
.]]4NQ2=P(bXRRDBJf;CK/<;5aO=A]3M&A1&M>Z-B6.GDaf.P.b8Y4RZbIKT^-J+
3W1,R.UgKN/R:TO,-VMW4&c3&+d.gH[(?,PBD:QdXAdb,[eTY45Yc-@\ZIQ6>#Da
JR&9/0QEf@GBWY-c3?=Pf^IP.F<#\>6TVA9+CLg6gD[/[F6EXPD?JGOQ4<E+8E[0
#2:U.a,0<CW;WDCg42F4deZ\;AS&,B#D,);SQ4\?B,PEeg?R5NT_J)9K5LUB?ECA
Gc&,QgZK3<Rd2=;Ybba:MP,8B_-FPS-J:fQ,=^&^Wbb\[J616\W>OFW[S,;/EcWO
aO9QGY5J#,cSY22YRUbX,4Wd1c4fd)PY_-^/>b#ONfHJM/58EP6Nd9XS#?WL]LYE
ceA<^_GdffQYBfZV&TS_Y1KV=?H(0?cVFC<#WBH6(d<7e]?Y]0gcAJb)]a90]P8?
Y;XOTV,996TOX250N^<@A3;KO&G^2(HR&^dbR3YRg=PgeM.JSD,b#HF@CeadYNNM
eeVZb7?c7KY/I&&E\.7O/V)=5.E60,2SUY//@Y;,=Z;+XdW)?@fC/Q]fS5KHJ+A4
HQJBAdPQTCfgJ\,SAf,)/BHDe)GbC6<<A_3AY_BV=0-FSH?=L6O@YQ@f.?^>CHdK
=7PFK^BQ.d+@gE.?_?LBU-O0WKJ\CNUC,HO=)C_P;J##JPacD>^(_gB-QJ>I<9=8
JGPaKYT3@?8=F(XJVc9D?/NF<^S#J)X00FFHR2LbN<8,C\<@Z.AaO?J?\7UVHcU(
17RYD?)Gf47Td[NEV(\Ac.@_JBgSXCSg]PZ)LK+G&ANPX3UQ5XK3(_c#bWVNbd:Z
b0.?g64L<_XFEa)CS[\?JMS/cY;ILH4Y[f<RF+V2^,1D3SSKa\E??dR8&O82,HKI
[\M;NI7UWYgC4YD0D4cg:NU1LIZH?e2HI<231UbaP(dcZYeY]T753Yc,[@=-f_c7
MN88\eY0g0J.BOf^eBX9(7Y<f0DI@E_WF?)CS&^J3X043c+=?AU&8@<9BA/.&aHS
ZRa9bK<gf?2N5U;PHO@DR/M95M27O#OQFNIcRT<F(+LCEg92K#R6&AcP@=?==-_B
DH+3d9=-b=[.EOMV#H?:XJ1/Z<IUWSb.[2><ME24H7GJUaceU6J,FM&GDOTG]f(Y
BHaSe+EV=64B_:C./4VNZYe]=.RbM(F4\<^V:1&b=SUAOg;]LQbXK,;b(O8MKR[B
7X89P]ZgD\SAdC6B8P,\/KU&,L1@1UUW2gCgXVDSf-MF,)ceSHLWL+#WBLC#.G<,
YFPAXJ&6AY-DETRI#KO+&=g.EA5;8Z7?(ZXU5RH,7J1X+LN-JgBG[6E>)-N1P;09
OcA>8G[V;8_HRD>?2,Y+gaI9_g:(89cYTTRE=<[Vf75P&(,-H#NMM73(gWSUOFQe
FJ6S):L8#QeSg3A+&4>@NW/:V\W&3+CVdKSW7--Y?ES=63\4G9dJ4>CKZ\UPJ8]W
LUC,-Y)g;J4,VC)@DJL^Q-.+bG[4WY[JYCAb&9#LHPV.1cW)b80b76),TXb[RTFW
YS_S0c-@Q<>86A\cdWRPK//JE?Jf&abAI-3d3MH_?]@,.Y53LgX<?&YSPNc=(EM:
-8-@bV@/,F\YAdbU2OEa42Oc=b:K6I6&7J4,g^14YG&,+(_C.aJa70e2CV<^CWFQ
6&2fBZ1+;42Z6^.[627WO:I07aV/e-f;9FGgA<V^IB].X&TdcedH^HUe2K8Ag:aG
4/Q>Y/&N#^SIcX2&_KYM2NT[XE)H?F3NFa#Cf_aPXHZNf+;gc;>N#KZ.G<)&Vc5e
W5]^Cb-94TdZaZ4XYE>4,53GfSNJ(0)XSY+Ye_LA&g)A=/+@>SR:60,3MK7F@;>(
9,,O8Q)ERZAdR+S?X-afNH=43:7:6W;Y:1KJC_5,O1<fVY?LN--=J1BT7?L_NTc,
cE,fO?PIR.M_-28eH\0)[0G+IU6+TYY0d[K1bJB@bB:>SG4E-3H7@>fY#P_2=I?+
AXB=E]@.g(bSO=N@fI3UW&^)R449[HD.1eNV?/d)be#?+-=/3MXQNHeQ+H?]>f:[
0NO_NM_^X24e2<L,1>,(T<T.e2e)Na-/(E:X;-AB\ZZJfS][.;E;d8c4L4U5f\>I
3+&,07P\fS=\Q<FgWF_#8HH(MBZ.g+7C9(02gISZ.YK]32JPe;>O7M)6ZOUZ5Q7L
)H+/O-5IH1c82OZC:4DQY,:4f-#9;\2Hf&^D,QH6H:>c2.H1&)GGMGJWG2[bPVU1
;F2G>X-VD^&72aKS<aRd.XKHfeWgW]]&O);..07OSbeNJ[Q\Z7VNF(/g)3d2>@gL
d6gKSHWb+DQRKCW4)Wea8A<]<(:eV<OH69GSN@4<G/O&VH\]6ALMX#EXW+<FDK/2
O;LW351XagaW#&/MCVb[T>6]KCYAPKZeKHYXJaAR;Mg^Z/TTB<>-97NH.fHXZVG4
(JWOBF8#O#[L=T08G^,)53IfbHQ]#IQT)c@@5XSHZgDg;Q^PcY?4ES02FE+C\A-D
3H6@?TgfY>FJ5GKHHSL/e[55Ac(<][^FZNY9<5eO4B:2+1E?5F7?fSC^eS=cdC;J
CbV(,L^2?F=Rc_S/#2YP-F=V(/[+JdWg#V;W_UPU(&=&VR_E2(WL0]4H\O2KcRQf
g#J]F2DX@-A7DOI:dbDLSMe7PFaI+)BC:UOB?Eg#P1K<).J/S80EBLSO5,;X+:[M
5?B\]ff7)K@Y&HW#D0XMgZc[TE#:V>6[W(bP1ec>5.R+g@>:9MecZ9H>OKBLa4/T
_RNNDFgOJHL@KPY;?.D+QUa,N\C[acLV)=X_K>BFKcCJU_&;=W#7SA+1EObG9O8f
U#OS;>>UDXOLd-42BJe8/,[]6)C9H\;0,J7R8;FC4UZ=TLVM0;cccST0a;0ba6G.
^8Ag=]M/P4@^Y\Q[W)]_#a,C9(HYf[FJd,dd5+W7E]>TTf^Ff&6;^TGMdc>9O,J3
&Aa\ae=1PA@UI>O2IU8<=.FF,-NdDDD@?A92PS7^>NEJBPdQ98B_W_]e:BIO054G
7Q7A<_]/0<F>FfUO_5HJRB^&A6Df#VU<1+NG)&H[KANU]09,<TYUd+eK>SJZ,a[Q
O3T>/^@G.FK4GWSa_D+8e>,V:S36:eRY[Ne_e>bCXPb.MEU>#JJLUX1[RLAdNIE)
@]VQ8:N3JCKX)0@]=d#<@&@4Xb5CAea5H7F)Rf6eOdT^NV4LfE-MT?U<^\/H.-H:
61PfB;<f)]f?cX(d1V=#5Xc3M.3J_N00?\Y77A[[8dY8HYBGW&J:&bfbd5?77B(C
VM8=:c8T)#YaXbLILbXGIaE3E;])1(Q6V>05-e7#ISWY&IH>52=d)WG@cQ5G8[Le
aZOZ(4Le55RBaO?L?-F20WI^cKVSR.6Y##G:V.^SY.[C)]bD7LeF4,e/gc>TP>UJ
[?@[e6WO3Q_bYe/+]11.?2Te&+RY6fR/G?67Ca1/LfGR3cG@/L]LHcE9:HP4e<cC
cLIHX#TE39CEK#N;]5C(TC+dRS10I<K-U6PGJQ;4B]ZIJ7BL9D(Z5,X2(U]3N(Z,
f1UL(8dYLc1g1GV4WcgM-Q7gaD]V7F97LeOV(e7U[8MV+XeP-XY&DC4NdB)7:><8
37\W7^J&Ze7+fa7gCddH/[\EZ,_1XDH1JF++B7^:N4;\(X(b(6Ybg.U1c9+F7(fI
a6W,:4ZN]99fSKF5SFF9).g?1GWMX2/fH&\D(K,7REJ6g]LR]6WUYZb&.M[2X7W=
Vc>1J2KMQ<#],<9bY,HOB9WR68Q-A<25<Q0IRBS9^>bRC><e)d<Ga[YHGEE9UQ:c
<I[b(-AY:QI4SAJ#TUe_Dfb)T3A;N.:KG75XgV)7CW1gE(K3E:(SV94J1=beT>Z=
IU+b\<bF-Z-;\Y6?G@I/NP[)+bB5+5SMHC7[+<14CgXe[E8ea,70V/V,(bX^DLLI
OV^;d]FM()Qc(->#(/X9]5K1OQ:OU9faG69).O:>#Xd_e=6GLSEd5ZWg>V91<\T=
,#[_DVDZ_3^fF<Z<e#_5c1=bL#ZP)53Z^;f5C6)NS-;(3?=W8,Y[(/WBG>H^Y04I
@f@9gF5-LS^B_)d/FZ=a40gMK\61Q\/A0)C]VINY3QcSC[;a2HE4Q-0gG=1ZW=cI
7dRa>.A<@U?^:^2/5])A7=\+1M==L,?//Q+D1R36Y#J^7AVTYfJW.P;fMQK[<7&2
\dI\VMaA=)adg)U9=&HV5_?CB7Bb0?UTFR1GP,N<K7_E\=RfJ+(C4ae1P5\#<N/+
=14O84;\K?AZPYXcf[=_FRF3YZ_9Cg:MIV9V.;Rb#YK2J7cX8<f&A^3><_7TNEKb
,M_3WS]J/3Q[\1B^C3(59Fcgf\V+)eD,&PB2JNQ(I,405F]5U14?V;dcKA=1M^R(
_^];.W?1a(EY:S8S=/O)@?9+6d;>MJbWHL#QJeObGe;+X?<>BSG+>/T27N6Kbecb
NYA0#B[YEF2_B1P,(Q)XBIGQDXCEc,+9<G)9+Z958Y32W4\;8Q+JC:35Z-6@RgXc
SK<SIY.<M<Hf^?,AHOEO1;QdLA3^/BR7,8)CVc/3P?H0QL/VDVg6OMf.AAJ97-Gc
6@g6@?YQ)8=YUEKcNc]0C\Y),B:#5N-c#F<1576fQ5X?cA[)RG[E3?XWM2RWfR\d
S>)]+X)FbfF-dV6;^E4IIgY9A>Ja?b[Ze,JEAQ+._@ZXf<FX[JNH2(8;_22]7aUY
_,?596[3b-XKIFbbQDaH8g^PU</V5aFeNO.92+>QNPTJE3+N.F<RBS.TSCaY?]+W
M<U[70a17,AK<D(0@X-WNO/aA1K#(DGH/7/@MfIR41SO]M+F<ZcFK,PVZL5=K_b<
[_PKR27(#[VbTSNP9#GH4e]+;I2^^MDTKg2,d<I8;P]\eOC&g;TV@7^^9->2W+D[
JHUY^KC_:E8H]VAP;9AVLgWTJIR2L=BVGY(2AG,QD6IPR3F-d0Y[OUSQ9HQO1TRN
H2D,a(fU6bKegMF4K&EaH:;41>>N8Be-_P,71A>_[E?8W8:f+Kf)BB,JfL++^KR3
:\C1>O0FbW8<DA>-^Y</69TS6bUUL+E4]6SYD(YFbV\GUQHf65.O;A0_TaD8)KS+
I7M.,K>FSQf&7d#HEY&f8\ILN7J+/-fTY1E9;;HC)1=)QZ-9R/NHN0FZAfYbC\c3
I[G/<L:0O&>&_bQCR[BYf4]gW\<?\&-D?f/R<6&G=TIf][[fM==F3KIOSQb(,CN=
;dVAbDQ)^-Q7V5(E7c[+=5R;f=MYgVK+BE@[@8/fI5CVf:6;:2R;R(\DJZd\UI[P
:a2BGWEW/4#LN\2^SZ:2XX3-Y>(H7W]6g:Xc=GNT\&a.K5E5M+a8_fU;^F0IO+1U
Yd\M5?\]DdJGV\[eQ:43XLAeZb[AO)Fd+A>aV<c=&IB_(_W0Wg/7EG5d[052Uea.
G:FU\#=)B3(\Pc]?5)]VZKDOZP?J]WDW?4_DV/_=#2f#@0,V2U^[9bAKE&)Ob;A4
OF,I-QC[P,(L&E/^M(SPCNFDU90BS?JRVWCGP<6RXJP=/:2,#4S3P\UA:7dD-P33
/3T<_D=3G(_3;VN>833NNZ=/[cJ\Z/:&<>C2fU0J0\JL#YZVPgJ]P+P@-@NUA@R>
;>L7/E#3ZITbX8d,.B/J76K0g\BMJ2^IB\>RTPH@;>9M<K]XM]WD7(F?>.P@>@HD
D#O:TW>1(1&&3<<WT)N[5#Z?#\J#0b07;JM2X[P?9d/[#-d:./4XYcYF.)dFe0ab
=POHOA2,9,dWKbM>5-9E<>@d-8g=AGJ>6-Z3_]OQE-^)>3#I9^dXOID5;^?7c)b2
R_:Y.>J]0]^C/O;P9\TgFSZ59RZUHcP?5c#)Ud]<>&T^[<FI@#gB7D)\UQO-MeBf
#BHO1eAcHK[@,ZJN-BJ2+LeQC0)]SW&;Y[8,OCbQgU/UQJeU/e.\B<W(?:Z)PE+V
bb,2dRWKC/[L,c?g+.)A9VWR;C(0eS8?)=#.3.K3V,E34?YB?T+7.3)g34>L_GX-
a]8aZ8+_1L->&9LPIW#f:-c1d2C5@df\S[JNf^;CcC;P8:<K>2g\2--B;2Z_=Y/5
Le;:Kb[-\:7\e(1HJX>e?RL;,[VSX_?aA5(EZZO?G5O=GF;eOOIeMSe[LNcd/,/4
9G+&IVD&)#La[g@&Q=^1Z:d1ETN#fV\T#QDY82W8)J/@S#2^L5YJ@I=S@AQ4+>=X
I?JfJK&FQWHJGgNE4W-N^K=6WN6.H6WT&0K[d\H)U+J?0e@S9+?/0Q+C\W:_@=WV
7e5MIALD)K&UE&0UP)I77c&DZUN@Yb?]LC?#1+EEE/KC3Za]@bU^d#ZN+NSW=]T)
g8f-I?b=T[_)d&L=NK;fUe)0IOJd\Z11VW,bU>EG0Y8]cXU6_Y)E\^?EbL1:W6BE
#,P6QZfN1=T;AeP>-K&E?#fK9;f,QVH>TK2?8U](U7Le8b-<b)&E4AP;W91W[Y#K
HBY6XW?Y7]f;=ETbZe(U_F#c]>);c)Y5ZJLdK+T]bdN8<I2JEZSGPG#J4ZMHP+^G
e=VcDO9I]C]&F5e\^D@NL8I6aE8DHD+<7J8>KY]c5(=(J?;O5Ob==bDC9X_8+fIC
VG94ZY#IOdd(b<INE.H??\Nb1F\.b&+bdXH/1M^11&L4:\)#\YJb7479,;#FbHX@
]caS.MP&K=:0D+YUNdAK^L6?B7M-c6)JY0gJQRWM8UN?VKI81YIWf6K+G+RSCA>X
=[OReR8U(X73^N]W;;K9K0E\Qd@T+d&<-gT)P3-N)d+BYXGX\3a_]Lf<:,+-#5?F
FJN/SAGV.=D?N&_fWB\@M?\B+[6a:\T6eeLO?YfITX^YJf^NdaV,(=J^0[^PJ5T>
2TWU4_,:B6.5X_^Geb:)HV&-RD?;8c+V9PbQ>TObCd;J,+K_AW9U@/Ke2>Q]e?)?
A-1[AGLQX7(0FU=JaR(e9AV.6EG>./<eH]9N<:=-_1[&MWDMPAP37_GLP\FB#_Z=
WTK&7gB:][?)I3OO3C]^6.?>f1HYVE:WU3-,6?Z13HGNTA#?<Q+W=VDX/48d@L-,
DdJ()QNW6?[.KWbUJ9Te2:K(=cG]S,3;>4/Gc;&aOUCc];F=QK6,4\]X^I2=A)NX
BcQ>K\_PD5BA_UG#;1FJHY&UI#Va4M]_.AdaZ=+WUc[JWHEM^^SEH2?=J-,CAX1,
^F64b[(G9@IICQPYS7FQf^8FLS<XGT\.#FdJD5D>00)/XdC::d&Jbb47dBN?QWO?
c_MNUETSSbZC5Pc84R0N5>a4?3A74bKI6QI48OUQC_6PeO2MgH,1J4Q^;AeW(7ge
Ad&#_?XY59GWd/&cR#=_4B<(G-3X=L#VO>I@+Y46aWE326Z6cgCUg1bg9&76Rf2g
RWX[@>;E8QB_)T&DC4K?8:bae/>FH2H<(XIAS[64ZB.gTY0751.E?S+V2\M=DJFP
TDfa]ZcBaU0)Jf.cQ[5-U7B6H@a.2O(Tc-Nf\=:0>?=6W(##M2/H&Hd:YWZ5,?:a
>IUD]OV&TJI428ZX^ZLLdZ)VgP8B)^>A53YZ_K9IA[L)A[VF4/:Y61/X&P8H2LH0
cO0Z[N\#[5+9:_X[8J0+YKI<LTEA4Xa,]f-fOF;>3T.ZdO4<MG)X&;2M@.g76+A^
7LAVOg)^;Y,ZJ2cPM+eeS#I:Y1,(RGG-CXK>X]YFX99&ML-Z4)26_+/.UHc,g6B<
5662#;QX?WNEINaW5L+S[;:+3RQ.)29B\CFOAPeG(SC3HU#,[YbRb(_WG8H<,+JT
NQeKaabBY)>G:#_HJ,A[F]-S&#eFM#J;+<,A;e5e@B)Ngb>F7XK-,XcX5=D.gJ&)
LSVE<e4IWGO#PKgPC/Z2bG.]?bT3O:EDW)c-W-WH=+b?M.W-#><c,2ZI(/JHPEF+
>CQ]IU(aBe_eAXfY@)^J>(L?N3\I=7T44WO+Q+2VHN2X<#E-W1Te]_:-(\Q=&JKF
C?NCIXaV-a#I,8Ua9cMdDIb(QS4?0CC5A-/#J=9..F)c;.4K5-#\H=)+CR1FGR^&
ZEa5J<H\L&BJCfF@,PE/DV=7a;TaT=(baMM(/EC:6B>>,f[P><QC9[b&bN1^.2b+
0aCAceO^c=0]_Me30#BdNYW\<]_D(#MIFFX>#;B=:555IKA./4A9aMcL/>BW,:6P
?BK,f(c<1:ER0_#J0A@_9XD6Uf5>,QRa]J<A/5102LR6>cT4Q+@eY/#Q33T;^4S&
a4M4Z]K(]3/U4SFa7DD-=GQDR_8d,[G]bdHQYFQacefbV[=:>:_F,6Z6/:K]1FRf
P(=R=:SB\La5aI[WON&QL2c\Q[8-EB:AC6IB,c(_<b(@?M1g:KZ=Af\cQG];:-&:
1,]+H;LL?ARXA_9G8Y?-@.@,98?+ZRVMAb87I#\U^ZNI_ZNP6<O1G/32W,2Q[0BA
QM<;1gE2=029)O:#E\W@O56KED>dIO=RJFU+:R0MdB[45[X;,G[]1_^19O5/BD5]
&3X_gTL9LP3N6MSBAeJ=fYJLN2H50C17)NCYN@8]ad?>,&AVQ9&[B<=D<I.B98AK
>Md2GQEEQgc[.S@f^6/5C.MTNZB+,.5U2)1Qfa1LOS5]KRKSaI6dL_;,1K1RTaNJ
MX0Q1#7<D((?]?\0DXJGb>_A4G8FcKV]3^Bb6^X5Q#J](S=K3032>X\/6<g-FTQ7
FJZ/EbV07X.7eJE@CHPJ]Ud[8?ZP)T8X?2+E;BbQD)TY;WG:Ge;5[GNMZM)\KXG[
;F\?]d1>Hge3=NBM4+<ZDYZea&QE)HcR[1+gQ;3=N:1(\9,TH<KWH49)G6eGOC2\
F+3R9dJa:a&dK+H75>bf._5&D_Z0S@=H]NJ]B2RN-^WO8CZ#BCVZ&P3c@\[GIIG6
3R;b9F7NA:-VOY_S\75N8<HTNYFG(-2cUBM-T17>TFGNUPA5VLbGG>KBZb^+ad7F
IWZ6SXAT5/ZLCf@0dIPdE5bGILNM6O-Y?\Mf4HP#PNU=HT5C,d]9Q;WE#UIcf?gS
(CTF&7aTYaMY^7gc_UQ3/2;K;5<&_Ze4)Wbe_-b75Q>9.QDZd\\ee236EC]2b9Ad
#Q[c+(::(UFaF/>SPXU1NTRS+J/CQ1B#[WFI(Tg-@)GD88M:GW-0fWOB)D(ML;+K
2&7SY=6RFD<DXND]B4<1-G]JR2b#]cU<^]G.0[XL:9:=Me_eTJJ?eP.<5a^;3:a5
f16Q\+>@&N\NP>#2Yb@6K:Z/:Dd=3]&-[.SV_W#?/;)U((WcEb7C(>XB/e1.7c_(
7ENA<b;YV:3.P>RC+YA>21JR<[?N6<0)TA<4)<;VFLeOP8.dWSF;1]4KMQ0ME-#Q
#ED.OB\HY.C^[.c<_CPI5S<#8VVVOM#O@J)LHF+2QGP@Lc^&9CePb)QCY8@g=8X^
9db(M6TS,e@bc1+/B&&cYTZ=^HbZ+]FAeMTL\D[])(@bG;3/KRX[S6OV<N4:V6>T
+TUcJXR<&aeS+[,=4E9[S(LU/c1QO\ETUaI](N=92BF1gf7@cM\K6K;aJHf-\P7E
S)8,-Kb>4A+=Qc#@GP>Kfaa-?S4TL<=\7>R,-.OK41Aa0^G,.44a#>(ZH@:;_=G4
SNME.4N8b)V^eC/B</ZP(Db=OI)T.dJAEC<<fIQC>1^ZZA7SXaO^ZfKUY+7F-2=?
6X\d^d_H#,A>8SR-dGCVYIea16HO_(DAPNIb=-W+(S,\OD@:GF#E,CP0VZfXNJB8
V5V]_7T:X;JNGf[[DN4<0N^5IX19X&6e&IV:RC#ARTf)LY.AS<3CZGdR)[)DNV:Z
dG\3Ja0d@c<Z0#S^QYY9e[XM)B<-BFEJ#IVSFBdb;/CVUI3./)/g\c8Ia7LE5g-.
M;d(J]3?F#TQ7]^W5I[@WSLTKMf#0;fRU;O8RVG4J:VTOF=ID+\&[N@#@b)6R0^1
ZHb3#0A1_6cR@3?Z?OXBeN\c#1[?:]WbWbI#.@E/<SH;[49P-?VV?H)-aSe9K9M9
PaY98KfMV6Sd9bV2eSJ08E:6L_[&a<OaD&_RZAgBa26?,126)(ELWW(SDEgKVP8S
:LTRW<fQ1OV+?eXN;)f=.)c\g9EO4@3fT8-_+(If3Ib/eacHc,WY:a=Z_(KeV9XC
3V0dg2:W7Y)IF2g?gF?(:A+-aJM1WWI2@4HOVCPHb+B]9/2B<)Se]\5:(&&G@Q0Y
NH)#V=,+=C3)=c?.#,F6YKQMa<gGZ5CdNc(U:6@@KSUCRa^<-49RZ?c/ADW/I1>P
0g(IZDf6T;3;BG?JGC:+2V\XML?4#.<3?U^PR5c=CE#.@.PcYS#Z0>AN^Pf<X9;M
D_cYd/UCC@:Db8d)Z&L(KSF]M4LX75]LWN6:&F6QMOA=L<VAeB=7+T&[&YNO2HVZ
69&=PT+K.Y;(CI7a20gZa,U>]Q(bXfN9=CGdbLJHgUL86cWaSH#195eV/75AON&D
3[g6TTPdA<DbUZV,^Ca1Egf-8-GJ4a,I_f\=D3\e)==B=X),^Sb+)([<(>U6I[+G
1LQ^3LIAT9/^^S6)0cO,MP.UJP>W4<0#&X))F;-U6FPD0,D:X,Z4)2JT)R@&-2>0
UFag/AOPSDP8d.ARHZ1SBd<NTa03&^Sb>@[eU&fH7,#gGA#De5<Gg1aAeb?N>_S[
NN\COLB6b\T57]O#)6M^9.:#M7TY/CJ@0X]dgb28TMf7EA\2R4#F5Cb2EW^6Y0+>
RbVIe42T_<:4b?-Ac6#eY-OgCR<eV4HcCJd79R^IQ-2&[);>_(c-/D?3#J>d\DX#
&H&>,(\T&Q<8RA=\YEIe);C<.1f)XYd#=5ET4f4Q&KAOV[(a:H+,4_gg+-Og:Y)9
He;PG>8WdZ8^g1EL9/FBd&Z@X2cV@?BF,4A<3YWX6aD>:e>d7L&[ALcH3dZ+[gIC
-]f4MMW(;=/^1N=8(f3F#G5#3_&;&+9I7g@dPeIAKIDE:aPdGUPO6KD0_YCc_\eW
R=KH^1C17#d2C>:B2I?-T[I=WTOQXR4Fg_R99^+=1<g/=>8/<\U@J_V=1PJaKWI_
Y:\1gJ>S&2F)V5;62TJ:IdL9eAFX04R?)a>U=&>>^^NgX2=[&(+V/+WQ(fcVg/2f
HKCM\/_DQB32S6g0GbQO^XS<VHSQF[O+GB,4FG&_\2:F0Ag3VHFbRg7=YT/@/GgY
X(G6#WdT=\E(8#YESfEUJ#TNJP_UKJUFE=CFOYU.<&BfUVI(HLa>4--];F;[6OWg
988DJ]VT831>9Ya@IRJ^(I.HS)e;,cY+J)a<^55X#F-]UGObAQX5\3]WE/EH)8Gb
af+gPOdHgfFP2^bU/C7-8G/^:OK9B@\^]&gaRPd(>=A0=#G9?5+GN2U]&.(e4>\C
.dU#I6]][VB#^e5[MP_SNMDI\A9CL,YV)3>3&1B#e>-SID<79#d<X^+Z.WE[CD[.
U)4/O?f[&X]EBETJG/(CT,2bKP2(0(0XYX04\XbeY)C(]HLA)DgX-ICd]OSL1HHP
#SD>P<7<13S>]HJ7I0c/8F_L,dEQR7RP&eD[KV]1ZD+4U-SbB2N83XA]V2/GJd4)
21,:.FOO,Ybe+(#Y4bgHFL_)M?dZ?_#^B5^b=7ISf1b/S56?ROa224Pa4ES\A)RQ
J40+dU>NR_:Z<3LWgC?K6Uee?1YJNZG-5EJ1_VWJ,B)QHSH[0Mb&f6Eb\AV2R0@4
+_DZ+R<L>IO)R=)e^.J8TGG)X&F:Fe]WVHCP0=A0N[a1]E=9BP:WTSJ7#4W@aMN?
9G2=\<MG72=,Ad0LQDT?W9:&Wb3@;EM(PN]=EgE-K0JFG@9D&V<A0B2.KXDO#4)P
<L5Q.(5P8Z7DME1(\ZaS9=&W:-fbbYd(W6_FgDZ3bL0&53.T3D&<5WFTdIN/67S<
DM?AD41<_10O=@T+_VZC(TIRRP,/\L1H+dOJHF^&fL<\<19QX./A_E@77^Y:A;SO
QcFJF8F/6GAU9[5^2<I#RFJN][7V\^eQ<].UQKd=-AYT@(W:6P>3JXG5A[R]VK#2
[@WeWS8[Q/Ag7J^9dESe?+V],1/S-I&CMbVK?5.3B6]VD=OF2G4=I@Qe\(8K\[A[
ZZ8B\D>UTc>Q:MJP(75TIgW1b/_I\M0?SB-C\V/C^HMV1]ES84Y.FD:@__NX<gJH
GW/:@HAB,\#4d236JE?HF]?)6W0WXL.T9+@CS6&aU(3E8bcD<NZ36K(\]Ug1#UAI
-ZJ<5ZF1)/M,6/+JH&?U0MX2S>e3\:<9L8W3QC[F2N1#dYI(8;28[U_5-A&?dOU;
4B>E:]<>S@WALE4BUf8:dMGH9dfT^,@ZYX/XT+<-@@^EH];A+23?EFEfJ]2^BH(a
.BT#bT[F:\J4ZVA@g]#VOO#POcQM4XEP<(-Qd<.0/SMg]0)#DgDES^H_2e)a],-F
T^C#b+3)YN)G\W)Xe5?d<C.Q@\)f>C&@<3gV?Vgf2RUN#)ZUP;;I=_e:Y6HZK,H/
8ENX7HOdWC7<<?d1ZOL?&e9.H[&W<cX;M?X?V3(WCKNEaKWc.Zd=cXT9XV4O?&\e
^RTZ[3UA(BVK9+H?&D\@]0-[9a?YS2L(:W8_<eEf/?bEJ#PE_V33U^b),.,<b^2]
9Be\ZN/#Kf&f;FS-06dCIMMg>)QMb5\e#,?/(125P\?Dg]JI][_fW6(-?MZ@1R_d
7?WH#WI_6gdU72DDK6IA1(<@bUGgIMg85:NNd[bJ@d9D+E868386]-f-a_>9SReW
>LdP&ad&#BG7N#CQ^dcNQ71EHd=Z8-A:&_>=&YUD\2_0P<Og0KQCJc2)S;I&RX=:
NWX@bJ=#.4DbV8^N,bDJ3=SY-_\)7PPaTP84WM3#FffY<LV_e#57a^_,U=1;W1H0
bQ?0ScZ;S5YHEbXKJ#[)g2EV/W9U(2I2Y.A?/?:4KbB71?YY.OR#Z8e7[<95)#KY
GZ#g#SS.@J2)YQbGE?b@fdGZC+94ODELf8(b4L#e@G?Lf,Y0;C:&WD>3;e0GLG_a
,Z\7Mbc3-.,:U\GFSMP0F[1KY;;/_7Eb.b)[HI23G-&)4=9_a683R&Q@8J5H=@DX
(KT\/#^8g[@&8=[W@7[O9:\VC.g)1&_D8[GeGJGK2:):8L\YU=7L14?3N_4X9H_V
PXP2UN<:6K+GLB.OF,_,FZI1Qb6(<P/->@a5EA7\eK-?WS4U-Q<,/26=1F#=#PCc
3SDe9CCfIWC9#;g-Z577;Za>SPU9VDA/P4DJS-A3DcI.=f?C2QJW9&4\9I[=33Zd
a5.LaMDVegTE3XOZ6)AfQRN=^WDI7ee)ATWUg7f[)TAb?M?Y@LO\>\Y?<?HTCg<I
L^PO[5UMN_:AY7G1Q9OH37e.E(W[NV[]_S_6Ee=5:b9(;N&J])=SY[)9XWXKc8Rd
VI@\,390f>D?E9PA@U/:Aa3E1XOS[0>-Le3W23#W,If3OTbND+>Xb::)&>)AI]Yb
UE5@aO6_P4ZRc\BTdaN#V/+TZSJSN_;7.YcT^9Fc0;575(F.Q&+QFXba(g.ENWE\
LV95YeF+,98-d?303/g>f\C^A;XWR+g?b&_E?:OeN0#]fXIT6T0bADR&>(DT/NKR
VJCQECROb^T&RG1.XE1ZFXK8;[:G511Td&Q/eZfBG@2&TG@)Z5F/9+AE_b1-?_KH
7FfS8Z58SBDL1]E@UPX&TTF8^PJLPN[\SYPQ6DS4cIZ-?Q7b?5[M,,LVN>;W-f=3
E<GV<-H,>:,TX;e2gJACGb7ZE&:X/<XCP3)&&]5D1S<)0W\?TV]-UeN>C#=dV0EB
S@f6XH/bYB9:+d]&cBL2d3dD]7X2D:.DNU5ZZ3)aBZ_UePff1UY_1XV0I/_;Ee5_
IKL#WA8G(XN\/+gQM)Y,+SEYUV8Fc7XF@:40VZ2J>Q+RRN)9[3+e^FY#;S[MB;JM
K#(4;6LN[)9+C+&4eB2GH#)+Y>9OFG+T-9ab9Y^MG:ZG_Y8^OEga,)E8f>+57IQH
T<D2^-bX;:M0M<d@;?4]@ECFBN@c?-.?f-<7[(]2RKg84E.Wd?4@/+V>a^BbH-(Y
JVf@T7Ba#c2\5=+MCKcdbA/]:>Eb6))-,a^4O>IL]gdfU7G_0W2aPe1F;FfVI?c/
O_)S]8/;G#4+1+D.E42R7MWP+^ReWQW9EG2IN5Mf@:,=5Bg3a_-)g]#.961PN<TB
+.HP.P6F0F1T9F^F(:NVfRT/g5ICaHT@-8:f:4G.Pb)1SdSK,.=6I>JRQC,.VVf@
EPC##MQ@.7SeHILX\Y+H^&#2^13#6-,C7M@?<D)YY=;154G(T@Z<++6?KCcK/M93
SfTAO;<>R.7318T5&2+f80Y2O+5D-^?:+?34+UYJZ10+Y)MM1---=7L5L3;D1gSL
PgY6=<(?aEF_3V+7)cgKMJ^-OB:&fGY(()2c)c>ER0@SMJX8bB>+B2=N3W6_[b=R
<AIf>Y()fHZ[.#BDgK6DS?ZL-[5^b5R7CXb79OAOQc+3UF6VQMF?:A2QY.b4S7MR
.=O/DKL<GGPb4BRJEH./(a])VPIg2LGG:QT[K2Zf[])JSM(faB+C,+SbEXU[[<O@
&8X3BcM@aGOK)8V:TQ/NgFUe2,.@a[F60>4IHJd3d>7N&+X;Odb2-N;=_2S+6IRO
,=KP8RP/P;+[7.^^#=)2SH1:cP)<J&3=f1;<=EEVdFM,d5#=9IWMOU\#-2;CFfLT
b#UY,Fg4[bW_DTSH)^D5,e+CRT+VS^K18\EfCY^\;=^9fR2WWMVdHCV,>NBJ2^c^
<8dYOJI91gIM_90MH^g?J<#G1RXcS>QBC/]G=d6LcJU/LdO(/V45BSL(W2?>#)Cd
TK#8g_.16Ag/_7B]<:C73WJMAReGgP4-Bc539(5.5A:\/(WdTH;)HdD#;V9BEMac
+MO,1eRdNcO0G(ZI<\..GHa<:;V=<)/9(46EN,K&,J&#\<+.8.O.CdCV@JZ9V-&<
#gd:CO.Pc6a[_7W2?b;@-U)M[2@=XQI?TK=1(K<\I<_NRfO1C(SYc1#SW/EV1.+V
Zec.S4N4CZTJfg87JH1(=5Q:4;Ie[G:UV2c\D6P/>_.f\8=U\?/>?^^7E^G3>U;L
@YV_BcRZ3<0>6c(>E[7Y<:Ncg>BPG26S#:Q<7VaV(W)?Ke^?UJ,+&aEW:U&X-Qg.
#2[<>OQ44,:,1VVIA/@GJ2d29>EJ46@Q+c>aD/g<0/=Y._6MXW\4CHRedP8TC5g_
c>LdU(1(4>f&-@^(=3&TA]S1PRO4QJ+V)Zg[Z5)QXAOTe-7cace?&S2CGC(ATAO5
::ESROHI>_5Z8[MfTLGf7[)F@gQCA-[&27\8Q86d2N);2;H]\\Ge\d&QZNEB_YgI
M)Lg81<)ZUfg?6^SPXN,:d)gX2cT8@VFA8gJF[AcW/#8EN<[Z0^e.H_Se5fe)f&#
E<;dS.RL[bW10=c,PGWBX;\37RbR+J9HHcRe[GdRY2@@V?2T@R>67f3HP2_<L)&I
Y1I7F(D.@^B3[J7cTCU#7JG9f)T(5D-;KNHK1#Ac+dQM&H1OX:/,5aIdA)NC;F:6
/LDQ5JCT6EHe+P76C[dG3Lc)@=MY05U5O4dJ9-G9g2XY,Y-X=&ee_B11YONIC6&^
ggL[5@[8&ARL;a1Q\2Hc?PfU-Z?6fB]=8PCQS:Q:C/-WaB)5D_L,ZEbFG@@bJQYG
gY@Id<3@cV_]U7g.9Z01MN&=90fG0JKW4>48X_W^R.]^743,(4F[0^(OWY)J;+c<
d]T#DOC=#WVb>a2OCL@\PX;2Eb\d:OQbUN,<9B=94R3OD7(9;gHP0M:TC,Wg77ag
>5\C43H=^[7]=0:JF>gK>M+3&R0XI:+IOUGS;)1C=@[T&W?SVV#V2Vf[M-K;+;KI
A&\N[F34#XZfY-JA>c(EODg&CUg7>48<e^4-4/X6A6/Y+Jc0S@@Td^eIRU4I+&bJ
.R05H>b)(UNeYA9<<KV7Q(/aeHd[K)PTVD,AN3dgH(,3]#BYDB];&6+5#;>Y:^Ee
gbV._T;2C2e].8AM9#Zc6eO<^D.;P6+FXA<:ISZJ4(3c3U]b0:Y&<Z3BI\LABgFM
3(=K#7Z2,(ZL&<F,dM=b_\442G71LU&(b.L@DUIa9I=R>?+gZKKWIb,C10DL:ILO
059<@<3_Nc9]H3D9B5U)d=,DH]XO)>5=D0V4d-+--GO\cCb<-c]\;SK+N#6Z.=XB
)3TO+:RI28[?&_#H+@dHNVHW1E0PaF;aBB7^,+JQIOK0J,Zgbe)?C8[JY&6@Z1TH
:FQU(&bdEDL2E^ED@Z:A56;FaI8a)G@L8D-8O.^bFg)1E0S+;)f7#=?1\BF^Z&:V
(L)4e\P7E&Wd,:?OLc]2_E5C@X7\c:+\Q6d:T45S<c],_5WN,R/;]bTM57bP4&-E
.A4VGg\FL^\P#g?I#\2f#@B/>@]8VEd:?-=@g=/:)6^Oge7(#;c1L#-Yg;/8N?G;
_E^?BQBP-2-^^:,ZW\,4.MbB4WbH?-fcF8aHC5]6#Q47H1NZ3LJ;JRdHPcI&\&-&
+e1[6Y[0R-&#N3YB4.c;#0d4QS2>dU65g>G#KS:K0KE8D<)-FXK\3@V24&.R#FY&
>1Z@VY-?[))O;B6Xg2cD-O(&=d:T<2D/VE2;dbRfS&IDK;fR[+TP,1Rf2K.;FX?Z
c>cU)W.JUSQ.H>3?2A9gZ+C#RFWA#Z3f7\UBaIb#+&=8V0#D-:cAWg:0)JV[(CXO
e;3?g>\H-LA]5FSfNOX.3Z3(F6-.F_IO&[_Q7=6A13c>dR1<O=(NYb+GSKH/eK[7
Z:UR[2Kgg?59dO9d0,O+I3ULO?994>cXJB:8T5KcC<-&OfcS_^Rd:JUd@3H=)XVT
43;cgU6c\2aQ-A472Z=DeZ_;:\?b?I&Q>X8;0R[R3QY5S(fE4cWce>-4_3R=T7V3
WM6Aa?3&P?OLWXg7L5#]]M3>G@bOEJ7S5^>/=2]H[Y<@;88)H;9-gHS&gEgM:H#;
fT3OD+TbWNOAOOUCTZ-]H5d;f/G<-K2>^acZSY#[E>g-XZ_e#T8Y[K:Z0+A?J#b(
K+5F&#R+VScK]1TJD37[Z#C:>+-P>RJJ1+C#K/bQ0dJ+05Sg6T4>,<6JU@7FE-9<
e4W7PJ<bWS.[@GQWU/^Uc;)].fH:&YH\PUX<AEWQMUHS,LZa_:fa>dF\JDM\:GR<
>0M>BQD<X/Tc[P\2;I2O)@51S^]]]H9+[DO(T:=IKQ]C><N+-?]DNDgQ,DZ@:AMN
U,da0H1I&?CeIPa&bKR_H7(b3C>^G[XC\EF@\MeX&,7GS^6Y7<J6DWD3UD.bK4O5
91BbTe(7Mc@[B2=);><AF=cG.e[<P&MLcd9(?<2gF?<RCAa2L\8^J93,+<9,NS?&
E<#],_=(gO(6(LBZL>28BT&>@U+YX6.:Z9&WM50/L5J&?)AUODR\1[,(+V:I,5Z0
CVCf#//K)#)K<SP?6Q<VUJ2@)^_f5d-XbKSBb-/)XC+MCAGcbLX_@/X46@9X^T3;
\FEbP(EQg@ZC>:-7K3QZ7CfU&+#QcLZK5Q]94Qd<E]4^F[O(]N4U@M7:==BR=<Cc
-K?9>]FCZ[gR[C,]>=Zc-_XFPO(f1YJ\6CJ)UUb[=02;b@-JJ4==T<&<]GIZcX91
/?-0>IR95N[;,O2Td);Cf3E3@[d5F15fccZ)M-FTH?)ZXO&NI<F.A)RM\Q:^[Wdd
1N:I-;&JB&?;2F+T4a]8_HIG-(GW;V\M3eZM8=ETB7R#75OB@&>E0<5#94-BAYd.
0W?L=aYHRfVJM(>fMe..aHD-CW1\A4YIG9<@Q9HX>V&(=SOMO)2YV&)?)Q@g(@[I
ga.31JOaZ+8[,2QIRRJU_H,1+(+/QDPd[Y/58PPY4.X9>bd_M<bAbSZQ8fg[Q.gE
K^UM2O:fG^OY4L1CTd@@(D0M=R0C:a]_6AK,G-QfQgNII2Q:]33FZ\C1Q>e;YP-5
3>]JMY;JD_Y=P=AHY_O:YK._BA>&FN9.2CVC6#[JaV[4V\WW?I2Q?L2BcQ.,&ZWI
?DVbT=ONb5L_5eK0N1_400O)JW+1Tgdc>W#@e\SA16(5QMAa]NQ?3OFH?>c,C)EK
6^8A;^<EN[M.(]1VaS_b.0QW>G3d#bZ4?@Y7-JET<6F1#+ZB>??7S:\c#f@3^:2g
P4OJ3M6A8NL+03d;MHbC3L1)XI?[6J&VU2fL\E?&,a,fgS6f<_RHXSTF>04,G#HN
c>TYF5B_RQ[1PP>:,=Fb81/;OQ0:b/(WFSQ;F]^^g)(LXe_+#<8F@]\af([c.:_G
IO96>U[J7]O06PE>G/dCAB5T@Y)e0QLGf3+M;2S8&a9;.+?51[Ff3V(9:\DYRg]Z
WA0_FEE2Q&SEGLRS#7MeF[BM;;;dI,O7D.V,LX:LE]Z0^F4LVHZa0aM2+(?YOY2=
I=-95U6Bc3MP>c0)fe>_1M#/C57<4YcD7.Q)M1AGf;J)YE@IB)[Q[A]4&3,:U2CS
CT;c=Xf::f^FeO=M:6(Y?:c.BeQ(b04f]6HA<2\/C.4+c6[-R)9SC:gD^Q3B..J0
:_S6<QK?\cD-JWB<YT#FOIE#:5YYZLg_>9f1->K8]3fa\K.QBc_7b><F)NO:T\Q0
^J@KCE-bc(CcQJL(e6:34BBg.L2RUSePcBJU)+#^5-E0CRM,K3>7(b3NY_L)R_WU
U]5?L3)>;KI:/f16\T0>GQ-_2e_9=QR]8\#b\;JeQ:,)K[0KJ5:7;@0g[NASP9_1
b#Zb\^UY^g_eW86M3f6VN:S.J#R_6E0cB1/HMX5PM@gEB,YgU6F06P6,?1QC03K:
bY71)9]&A10N@OD2#OS=S+N&2F.<e[5:YBDP5dR8?^&He?VgbUJ_Ge28716CS=(/
QN,XNgc9#]IU]Z#[G5]M:#Id.g:P<G#]F:##X:]+EW+POF>bcC>8-][^\@+Y:1QI
;dS-dS7]#f_J)/ML.L8A]PCbFUNBN+49RFOTM:]9)TU&YVOEAZ;QIJ3_A40VE\+3
3.BC^7g+SBS86+4Z[(S8feYSGXC>+B\.IB1MYOONbW):c\g<>O@WB<M>H+cKXM:.
H.1FX&&G/\93=/:S7B5LTbPB?IAE?gT?8E&FTK\b7Q9^CH0?.)N1C:2QVTD<g-&Z
G+^K+DAKa>a^=<BP@NaGaE&-JQLZ&IZ\ZUX)V#CbcVPBC\#MIS(Q&ERQ3\4CQ4gC
V,g:Z-LTII&gY5UYIfX:Kc>cE:A6L19E+e);&)6?G9f)->/NK^KK<VHI:D[Y(gMH
T<;#X8d4:38,B6F76&7Zf0:O6J[M5)&+M^a2\EU@C?51I1&(><R\>L8Vg+03(?3F
Hfb9bX98e2M=0BPN.,<D.OZSbVfW#OSS,B)P01+7T;J,6T7+@9/8gBYZ^SaZK/Wg
)Jg+F8,_(aK5\-2&ecF>JJ\\_\-3?V.RGAN2&YG+g,cTN3]2_c<7DO+?Q)N)B<V(
>?X8Y3Ia-(H]QG21:JTMRMbe+=b=_V0_M]HEJd]9/V4MN#Ga#Mb]>[PgR=.YZZ72
f:\H#94)\-gCN]7UVZ.Y6Q@fNK7Gd#a]9+_@gNP7O6#ZYD4b)M8L3f/W)J+?1&eU
(J6,R]=]Zfe:bY.0E[\QcM.64E(,227@V^#Ue/2/:/F-5@(3PS3WLB[B9(ETMMUS
ET^HI&XZ_fL/6;?9=ZbFS;4YLeMHbETL5+gE1U/B4626SE\O7ECA4:EY0,gO.I@[
0H>7Ldge>ICZ\\TO0D?0e=I5RH7C[HP5.)IB/-H?J/T]_8LV30:DRCCCa>3]I<_N
F5YAgNR.e074_F24Q)U4GdS9WL>[RX_<c?Hg6dW_:9+O&HaceZ=^=0Kd_b.edZ[c
DG#UNdg-HAd9+Q?:#91U\>Q7<>b6>.BP7?]U73:FOScc\7SKT7UV(TVO7Sd/KG4e
JSE4W:2I^][0,W78+0L_1cH_R0;N]0O2OSB^,Y@)5:KYE#3A0HH46c5B:/A:X_AT
9EW?C<H3AS323EaA1<Lf2TU,@-Y[1AcZN+=#CA14B?V7DYRV0bO_K=J@GCY[&8SU
?;7c=3eR3>,bI,2e^WZ[dX>[WA1,+Y(68W+Y8:/dP=dIdCH_TI+@SXeM<F9SE49.
&b>U.<P1.I=eDg[EBE,2.C5H^2;6F:?,7MDN.+IcPLI4+:Y1EJb@?\,PYS\IGW>f
6H[SZ7Y6]S=4W^,H.A4;ZIZ#f4<T02)fK+b@VG6>dB+96T6]<0cc@YI__20R1KD3
Q4G/TJd5cS/=g;@.0e4+>@P_=20a^B(^JB-,VGQBNJAf@KQI53,28\CF(\HA,JTU
NEQ.d(W?RTAb&bLDSfQ?Pd(T3b(@=bVdCTU0S-bLS)=^WJIG&&@d)-&.ONS-a6S^
dB809XRe@#^e+@G[A;4&Eb033_39\5.Q;Xc>W0VJW:CC9<WD)C0fa@fa6&HHFRYJ
\HX3De9J:e1>bVT0X1XB@XE?ea@b]FZ:G?SFf=KX&RN79_@bD.D?#O<)I[#G_aX7
(_OJ,>)+dD9bHIT,Q42]C[>^LKBU>):VR]/7W&I-O-7E\&WA^EbCA^K1LWV-KX3X
-.#1J_<H+cV?F[:;?9)SZHO?\gf7]1>04ER>#BADH><V0[O^?&L78U5\>NX;^RRf
L2@RdO6Z3SX#1^.Me#4+FLB@5)58<T2HHc+Rg-PB>M=;AA,>&]B1Q.[)Z/5\/<GG
8U4ZG8[We.E8L1Xc]ZB\;303@<gQ\UQODUS>T7,N#G)=UbdD]6@1cYf)ATSd;QA?
PG_B[1XJ2@.H^[4<3S?=G_A5@JQS9\SHV)B>4KL<=(Ng76e]Je3N.Xg907/?LHfI
?5>&dX)=771W2gg,,(-/\V.=649V8afY&3)bHA&,7=V0>3]AF#ULf;F;Y(XN16.Y
ODPH6Oa9QGaX0RFb4X)\-E@^cKM8P;SH^W4,<12L4V3573YY[D;XPMNc6).Ca70U
KY_GM,7=gN>(DMcgd,d9AJZB^UaM=L?Sb5Ec4D((5;XH>CC?AQc]QNAMQ?eD@YRW
S@Hd4Y)/]4TXS/J<3^SFXZW<?fPZW,MJIK-S99PV#_Ca_U>2\O>eOIBEUF424UQP
OHO:gVI8JdU8FD^4d#A#S,XV/?E-L#Y(Z,ZgL-g4U#^\V2\:FLeE(>3N:5&0&-a(
=PWJ+(I#B[]O9RXX)1HPM5dOa=BT9\EcbHRC&U@OL#-9>G>VAadO@E(8<IU/0T4A
_f2efZ^-S:O7?Ie6BPd4f1:HRX9C50^^FPF9cGWQA/LgSI(LAC-3VP:E0cJ:6ZJP
UaV)VM124L3E:Y+\66&S-.eZ;?;,N69+aS>[2];T4U?^0H;K,+/W>^=L/^\8-fPb
?95XM4&#>>63R>749)W)9X0Z\aBS8[3.C<\N-]Y?APg^:fOgeC8N1&\1.e?CK<g6
R445D93Yc_)_a3E^Q#,>Mc\d^BU]fDE+JMJ8fG=T3@HTZ^===7[4#K+c<<)g95,-
9P,JUEFCMdR9-DLIYVb8Z;TGGB2A>1b>A@:4GG3JWY^<O#ffY=--OU>]VSd5U?ge
8V5fT0DSC_R_+GeaO0c=A)(Z/PJ40G:0NN)N1_,[BXA=,M4N\F)L,,,L(Ib^P530
BVcFRU4[KSC2,0/K,?4E9#:F:DL);2:aXN2)2_.W36W??C<JVG:f;CdA\0FQFF;S
bCP\bd&gfL;;JbA+Q-EB3eF,FP3Q]E_(;IUP7Jd:UP44-I3SIYW:W(9L^&6KU9,H
_Kgf7F\,5;/Z=G90XP@4;)dZPYN,U5PP5Ad>X>V1,/LFB=bG<OE9TS@8Q6dS7=\U
eMXb(W<dY.C_J&-Zb)P5]A/:#Y#;NN?,SZ\YFg74PI?3=70\4TcHN2Fe8;VP8K,d
;;\()CN^UCP-(:WG,/J+Pcc_1:cDNF=S#D;(K-:U=J.H6O@8g,7GD/G[cg)305D_
FS3P2/GK-YGaUOcD8J3=1SD;#9FTC1b9>T0c6D&@dNUcge<B+1<3;]YA,+MZEVRR
SM^.&1H0__5Fb)RQ(&Jd[T<E[&?aK#=BL=N]PbJJ0SL<g?X3>bAYA;D2OQfM0eVf
E7MIYN;ACcbOX,Q5Ug\-^+UVAbR0J-(]X&O6P8HFZ7<2&7^aR&)Od@<?Y(Q)eMd7
4g9-W9H_D0GM.EPEJ]d]V60ZaOcGd^V=Va=K_fWGPe#A<1c:1)OUJST;;C-J;WJ\
&NMG,Ec@&&gXgMaRPO/^aPS=)I[Od5;V1RfLFQ4\9KBFX=b/R2L9HP144a93.2O,
4,GCf&TY0#B8(R_=W20YeO2Z;K+A3H6V<&(K=AGMUSK,gD^N<=]2fZ7[C(NO.I(P
2W53e46Bb]6eGBX:CY+@=g0IFG#g00,e@V9=B@RCa:;+>6UbV)Q-AQe@;A&8<LL2
2SY8ZJNC@MNDf9V^@,96,L>]CRQ-:U6567THe#[738;\aUXRCO3,A8:\b(C@Qg(9
JM^Ee]]1.7<X,J.1C,_Qdc_VAKPM/8^9:#]&ZM-&H87R]I#QI>@=K-B6(FV-X#@:
5,I63G\X-PDGY=EQDTYPD)B63BZ/7BNGOLN.KH_6#0\+Y(B(W>D&@-ZD;JMB)0Hg
JN;g4fLDXa2-UZG=7a4\K,XMf-70P2g/0+a]-[0^_@_]MRLFG_^-XEK#0S#^?\.5
=X<f])TM5H:.g2QG3LD6RB_0?d(d(C>9Z^K8Oe@BL49XaZ3L_ODCBKE7b\)KFaT/
9bZ6TSC]:4IWc88\4db0eT9Gc]f#b>9+UKBDf)2eNC+<>S>2:Y]BA:_/NJde=eE+
6GDQ/dO;/0GB74g38gFK/]1=OAf9SK&Z<_6100KBe0/Vaf=4(+3CgR459HQ(X@63
1O5KEH,FW&0_Jf59g,WaJdFH#cZ-TYc0&eLSU,U]M0g?eT\1a]7)c,+(acW2baE#
F&S0O/OaO6(>8.[1KLOZXG(V1WD10_,d\BXeNa[Bb_A^7T59e431W0JNWd7;-?F9
K7aV+1@GTG7b;@H=_ASALL(>Xa+SWdLSa6f-2@(NXfYB4RRS_eTKW-2OL6/<O\1c
@FW[8aVa=\D5WH4VgcAT>(?aSQ4-0P7E-c(?@5EM8>XDN0/QEI5E_R?7X7-RS:60
;,dg7<BGN0eY/M</f7GY/E>&LA-@Le<a8ab4Z7:1Gd4d1FCWd5J-g&8@g9M#H(?-
_Fdd3>;bT,Z29.H[:BD:\PN>HW)G#LJ;ZZB(KZ?-N5QMQ-\PF5I#Ag8Q3fG-W:?U
D<T_F_<[TVd68U21)G,aFYC3LbdNRT4gaE#/2DRePcV=0Y6L.LM([>RS:V+eH.S3
N-Z>;[M7Kd>.P;8@869ZdgLXWf&#;T<dbI51;Yg0+A[4Y=JI+=TJHfM,XL2S[E+H
.e#Z4J_,/]d;18\40QX1CfW\SDK/PL0YCN7]?bV^?0BFQ99fWC#-GBgL(&PL77<U
KCX:[X&NV7DEXFBeJB=++BfI&.,F1GJ3gF&43dbAE41c:]G69<I3W5B1dG,(e#J3
2FF2#4b/+@5M7Xgag]RBJ07.?,&Uf&XW73I-?<>XH+-D<0L_A.BTX7Q&Qa?^Rd4_
G9)<KAae)RfOZ?SeG)16LK^H9S1N7W/9SX/?8M]RF.Sb:_KR(2DC26J)^>T5GQZ+
X4c4(Q:ZKXUbTYIN3]7SZHL4W;6/40b:GIB70MI=^B7<<2\KZg&?[gI)>#Z/1&ZG
M6/-Ha26@3+4&1C^E65C\^8\##B<8.KFLTR\_>1b/ZDWCZSBTHYT>[<=K-0aLJ_+
EbZ\f;(4H_58@V:O1Y7V9TX5_E/(g73aZ4gVGfCC5d8?CA8G(^AVGQ5_.:We/;A0
.,9GG3A5dN41GeY_J:,GEE0LcW7JSKd3>3E=F<L.@)E+=A;gUYe/cGYY1J<L6beU
gfE\;K5]g,E>(A;.2N[bH@-Y0L2WfIF@RI4PM2&GYQaWENLRDM993W=[(MWg;R[4
Z.c_S81U]?>;==d:4Y4fJ;7G,8(VMQ[2dO[fFJ&Ta-;9Q48:V&(a12@YD,Hg(@eC
R2L4OG7GINM\?97=#PcVBD@)C8KB2T-:J^fMIfK/Y#fPTY^,477SLBcg=eBNc.OC
A+#;f8>gLM(LbM#DE[O#:dacY/<B;KF]\G(;QgeMP(L),1(R^_+N(8gS9(2.Z.,:
7O-a3SIN#N@4BacEaR\_0>T5P9^g#Q]G?eW1USJDE+FC];aTTX7I99-@J-?R>J&>
E+ZcB\HbM5:0JPDEXeXdbcTAI#G&V3XXGD.Ya7LTH^E0&)df845ddJ81H0/&#94@
LMB65_@\VSO.SHDB3#G+dE6N]X&A.[P5Da^1S7ebGP@@)86-IM#V95OR3?78C3X.
CaJa4IGc[fPC6C^^J&eOB,IE.D.R+?58[9X@fXA5KJdSGW#>@a#CGf;cJ(HZU>P+
JH./e@>GGRbOCTeFA,SNT/F[R_\G+X?-EO@S,:@XS<&bTGXDFd_>AQ3V0&1J?WY0
bF.VZ>>>9fKH?FU83Z.K>+H8SS,-7?7-RUT=QaU6fC4-LJ>\S.T0_QSQHUU<HBS1
[ZBL4A+bW3/#9T\7JP2gcUXg]?R=VA3X;f342<K>Y098UI0+J;LR[_8,]QMM\58)
[L+K#gcc9O3?N/M<fC6N_Pe]VYS;^cNfOMREQDbB4SR&^@(/?FDJ/RM+,@<Ge0BN
J>9#9+RZ@U=\@cAa1R)+8RYG57SY<YM?ZWSK\<YU./1J8&>:ce\HW&Y[)SdH\6LC
B).]JXNC\WgG)SO^F_HX23H/HIQAC<KFad<HfINfA9Q.@45Bf:Bc.5W3&HS=U&HT
Z\#A6_)<GBgP-DN?>A(#>Y=d_3/a)cRBR@eXY7,ACKV8?Fg-R#Bc,=7YG^US/YbP
3-WKJ>M&=_4]>XVGY7RWSL?[3_#D8=JL5AX9+53]#I=Z(_LbeM^T[7c+Q:R,U]LK
S2e;UY2&M4AHABQ<dPcc&cRbUg6>IA4(.7#XVb=8c<^7Q/2EPODe8f;TNKRa)Sf=
.1[W++Y&XN]aeV&@B:IM&YU_cJQTC<e&B\@F#K3e)C9@@2FZPDE,0HRSAOYgI/13
]S6:_/JSMHB7Qa=.Q0gDb.e:XGbbCDC(=0gB0?,)JDW,0V?/2/MKbG+-SZ[BQC)3
>K_+X=VPN7D=OJdaKTfe29Ig7b9QW_EAFJE;5&4.UMR,K/f]I_5IG&FE959)aCeW
_cXOFBVX\ZNWg7Qb.XML-Q,-];b_d2\\==aWbfUETfXJT_&+))19C00XC\2)b83?
/-;HS-TaG,2L,7;(SCSOaZEB8b<5\f)_=J3WM#0,)X7gQ?BOR2L[U[_P&6#(U+/e
c6Y2DB1TRSBU1G9+:Ig6Tc(9I\Ic&T?]=;9MN?L@VaYMaITR(L0&Bcf=MDQXHV2O
KAS&(Ff9Eg)U,^6[A?(9&31)a,@@E(B4SFAEEDZ;MJgJ0Zb0R6N8630M-#9HbAC#
2F9+PGJQ:9f@^Q/DXd+8(M?&;K15T-]8V:@8.9N[4BX.H]\8DO/-17gSB8+3MGU8
S0VUR=D8YH.J.J;61,[+,>T=HaI;F.E;^a/O\65ZB^629A)4c&M-F[eC]g:XN@->
41/G0JPY[R#30HM]FH55LH70IF8G3b[P@Kg)D:dB;H/R66.d5&;e^bXPO&f<5C.N
Ff/CUT)S>\E9PMgS53+9VWbVR0SI;EF8cb\_P;DD76(A(2?^T_T4;ZST05XBd[<S
I^ZN4_8MKP8H5c9ZW41_MB/2b3Mf[UC7X40L?0NHO/5+Z811?3aN;1NLG@H-.;Ee
0K;XT_-Vc0]-E>)TNS00]HB,ALJ.[OQ_YV:HJJ65IB59M8\8UN_K-P,C3=81QOZ>
]KYSZ[)60<VF)>8]^W\OT7^1Z[1]\g^UB[[8PHdWTLF:_:B:5_+Z#SE3dE1gG<\+
G]#HY9(V/NQH.#AY)b@8Y4e<4RT:I#dTL2a->faBAHU&Z0?NFIZb;Z=K89M36Y#K
J2ZIC]VFEQ?6dBWFa3b<,GI6H4b3/U2LT8.4VR<5[NKce5U,XN<c.)TP4cA])Kc+
[L9&X3<H=3+Q=B>6A7QP-=e]Q5]aQ(O4TR-821G=IK4Q=3)/J^HCP@WQIB0dKZbY
OaR_UQd6(Re?G.gY_gb-0?BY3VIL;<Dg\I7N)S0PM2^<&d8JK>Y/3Q@Ae68IK5=S
+V,D<)Oe-?\c[<=6Pb2e]Z+.e#K6G#Y3+gF58(&e5A0WU@S7A#1[AVaSA]0Mb45c
#-bAW@g/P+U<R.[a3H6f>/]_@bAN(.;D+_Z\S[K6HUG+]&AfWQOR.C^.B[ZPA4VP
2,;eL&(53I_C^PU=S8[e>ZRg1<IK84WKMBaR1HRWH5VB/I6I?6^M-+SY/aGSDRB,
3=EaF;ge+#+VWfZ83C3_A0V];3D]aM-GS;;Z7445d@XV0==g^WOMQ0c;2U1FL\4Z
WQCRZPN7FeJa2?N7Q-e&I[cY>V#OP3,)fC=.30<]UaL,=V7^;53)YY=PR5,[AJF5
K7SRB-=bA4g60=/g7:XOE2eP]22M5RgLWbODX;[(,HA0PR]PMI)-#:;b21@=9g#L
1P;NFdW=RFO#eOO[d.O<412LQ2Y3N&eJfI6-O_VZM&eHTHJ4?,239Z4D=J9Z2&HV
-L6bU@62.,V.E?20(>QYaNUa-#QV<ce?+-Y&L15&Db/X;1C:f61U@1S_/?1B>>=T
?HI@:L+R9KL_9&D1eB1DK17BcbV20GDe)YE[)J&J=LZ(f9^9gA(\K(4=R.6[O6ad
TW6=QfZ/eN^+HS4S8XLTbL/H_&=Hb4-S)4[RN)-JMQ)Oc1XBUUP&XM[/J9e95T:e
bX1]KcNXVSMHJPJ3HM/Od&]BEIVTB([b1839#Q+20/T&E(BDS;-3=6e9G[Q?4&_0
f(bbI9Y8]B=,])K-_VYVL849b5f:K^;L_1^.QUFFQI2K6TBKXD^19FCS7MZ&)U.B
6I39RCTad=RZf0+A=4N)XQ1ZPU7;:=NKN(c=FgdK_74?/[+Pg?<K517QIY]#[6>c
WB8-H_PgGM]AZ5DTDbSX7YZP2CX/^?:<(Q[A?#N5=N,YGdS9\bK/c2f0^P(:(=(S
/,W/RHK>6Y)9RO+4+K&0^Gb@2d34\S-XR(@Df,g#_<H6[0D-/bVO/;Y4V&1)EE+A
@X.5W-ES2JY0c41EbSaVRO071.98PgOT/DS5]2V@^C73BD:O/IWUEL=d-?5d=U#Y
R^Af[Z:YC.UT,,:6,HKUO]6+DB#0]TW+f=_B65O1PYH:5I=HBO5J2?ZeJdQ.LG9J
9O@,CAL&P@9)@QfZZRgE)I[B2N8Rg6b)L+Q(\#gP9GYfG5E]]@O^XC7gD5MPMK2R
TS(MI&S4.b\[_D]R2Mdd0P07C3APP]+&N@aTZ28QID@f\gT+Z_E:MM/gX9gF3++g
LAcS&E:Y#gH6[>-N7ca^0\30GUH_>g#U+cU.KB<>&.B:dZQ]Y.FYQ^;5SL@/_RG5
WZ8M?V->e4K5(Da_6RPgYPOg.?0B_.6WEag?\ge20G4H4&A^=4-;#Vdcg=dP:f[A
N&Of_P]g]FHN>^G?_2We5]/KP/TKNP3()g#6/6_gc>-9=.+LW9M7&Z_3d4:e7H6U
&^H0;GC1F?bH_DeO#.X#W:E9F+2W^N+#eU<5ZZPY+[B8<><<_TI0_^aF^(4RPY;N
K7RH(4;W13=4H61UKe=HCEfXQ1QWZ6Vcg<28(A)D8Ge18fb+4G2e7O-^@acd2P]6
NT)7PBFIa^?PJAgc?<5B@;58H@()H<Q#;-SCSA_):-I6UdJ>#7D&eAC;LLDKL_EM
5^[L9a6MF:4@3@-Z,fQ:/ZQg]D^&^Z[=a8KeV.WG00^eN=B,U;T-K>V&&8P([75G
89MQ.2L4Fg&9D^A,?Z]+\9LBJ-FE/)cR1WX1N_2?N36AQ9.42O&6EDeD)a-]GKGd
aE4X0AK4\R<_KHMV^603)23ES@1)K;10S:/TQbK\_Bc+^+RF7d-YJRc48,_SD0QM
RX:3SQ0W-#g@fQU\X_J=8I5D0<2]<dg[&A3a^K<>,;QFd)g8:a,7RJC0C&M93O,V
Sag\:.>H]=C72YX=M^2_<3-8d,Y#QEKXMIEGO5e#eW1WEIQ+7XH)^bG/L?/+G>F_
\FQQTg,6NJMBMO[,]2eS27=^>DT[N[]f;d(0Xa[Y<0A_7cKM_)8J#Q(ZX.8SL.PJ
&W#>^]<E>+/(/[KD,PRLRJ_<1f:RcPAKXfXg-7.\-XMJYK/F_3&,L7[HO76B?T75
DQT(a:]JM5<f+@Kg2YbGJ(eg6]N]eaM-&Fca]KND5+c#8,cIG=2&>]+WgEEd7?e8
Y9)F\IL1ELZ0.#Oe^G23FD+?bNSPA6F&LVFTE=PN2S56W7T^HY5,bF5#+d@,;.bJ
VaMPG]TNBSO:b2&U,6KIH1+;cJ.OF[H_<6fW#B@B+F9X16\.[UdedHOU]IJ?SWZI
?Wd0I^,B7YdU40AYVI1_YFU+5T(&bfW+.db@SGg.GBMXO+WS:#1BT_\A==\,+[3D
>?4c@0?E2gU>-fa@38eQAOR74C]DGO[_IbI7;[NfV\D]M6J_A4_)]G@VeVV&ZL0/
.\=dAGVPB&AfO]4Y)9#,B8CD+JYaZ<Q#CW5TLS#U(WL/6#5Q3K,M)^+.&WBf>.dD
+7)Z<Y5-UEP_:=L>28R^5<KgAB<3J^fZ8.^L[.^eQB[HGaFc,P1Y8_AaS1K0<#O\
M?=d6YOS0bfEBdG&0Ua:9cHU]]PU+T/3:d]b+dQD&C[cSAAe1Q.eY&>BEOH6X3YC
U.GT13NW.#618a9RR9RBJVPRPFGa/-g_2g]&R;\<RYGOY_F#cFcg\8<3OJ>33_?:
c>KD6U8&V5Ga,^-P2WCMJYY4f)-b[53Q_8@XVcVe_4P7L^I.P-NVg<6AI6.X8X.e
ZD;]1gI;9eB@[@=4IKFBe@7[2[0S):Ja)R/1QUZaOdWH.<6C-)SeK@]Ccfc7OZN4
01eJLOCG7?XDdDcQEN=acdbf95M[1HVc.I>YOOXZU3Z)BF,2F0[d>gZ&c_fbHPL5
VJ[9Q\=MFLHO\&/=\#9NJcSY_G6I[J?G>A=T?-@,^7db/Q]2]T2KL(0PDP&MA?6e
TS5YL6DbcL(WQMKCQ1BX#YHDW?ZUZSJ?c\cOZLCJ9<3O1S0@0^bO.TAF+6ccA[M]
_gL[7[@A^fZ8BU7B.-bY]M-6&YdGgfA,(E\L]1MaT6RM9Z3a[+_RdSAFA(e\=7Qc
#HHa1-84B<G2Bg#4a6+(9<8BA1AO2L1@B6BKK#Xa^Me9=aQ#?P42<HZ0\2aZ0d2Z
J26I/^60LA_a;.a<:.K&)87?Uc][;C=2NML_X02Lg?_<^BNPS(eD+XgF1c/(..dB
&B-WP6;ZP)Q8(24NJ<9-4([C^F5QKJ,1^7g7&b[XS1+(@\=<1=,F]3ERe&E=@91I
gea\d#0A0]6C4ba3#]Z#6bKOGF5/e+L#ZQQ6PP_UHd]ZNU_g+,C#_/0)Q^W]6LI>
)6947SWHaP5ReZbR(7F8eVESIB91Nb>I)cd(E9b.@X4[;8IHG))7#XI8_^+f]bK/
M@ed(.4d-]QEgO=.AM4)Y-<4Z@;5bG:>)N.2bGKQ4(eI_F=#(IFO,[Z[#[[Y<B0c
&]VF1@LBad2B.0D^bUSS7@A068-gc#;2.f2eV(05PDP4fLDLE-,@XUb52BE.2C[A
ERW3Z^fScR5)VL.DAb@#;UQ]3aWD:4K_<<J9>e<X<7>=CS([<B<ABeGgK9P]=KO(
F_-(KAV6K/1W&g>&8GQ:.H5_EP<L\;XD-W,IPc^P[f5D>)LR2B_QH23N#O4\5]YL
-@6_dATLTM;->6TVH8A4]eS&:EHd[D4<HT_<XU.&V(g1Ne)DWg63-5T;JgT<R;AG
:JbL4O2:gSddW;Sd&OPBG--@\BR&6MX8PeA;SJ[OWTgH?eR1DD<7W?R0c:5Y4@HC
6HW8?RN4f^#?fS;<&aO,PG[X7?<K38&HXBC(Rc<\0G9;<89I-<MU@+#HPY@=-Z1D
KbIQ:MLIBgRVNFSUF9eY9XVXOU9-b-L0PW8^Da3^N>:WfRDS>OU6Z[PI^NF<YC1J
J0RN(e5fDSO(\#/beKGdC)6QN:g,9R1\NKD<Ya=C]g1c3Q>U-7&DdM+WLL@==d:R
==Q1<KI0V\FK#QFD@\P87L5e)U;U:)_H8_(eGLf.1#cda<?-F\K?XY9V.26]^N4;
1._L-e3^C8W_T7WM[<)fLJ-94fBe0.2f7/[H4VAO4J3=SSU?K<777K1ZaB7)]M_P
(DDW9P9X@1O)L(NcU?c\=:T[IGZF\S?CE6_<b=UbbUQ]CcDW2G_VgId-=S2HY3Og
2LbG&.SQ3DA<E_dP3)XMAgXgM=(G^+&A816H<OR8ZQ\_.:3ZLP;77cRSHEM^M@]O
=X:]<?-bZ5W[G_<#)1aUd\ZW?-?Rca5Q2KEEB^YQ?CH/.e-f^\ZU=?EB.&H42WU-
Ic-fQKR^4=Ae?=<KU30accZ-)_TT\4b]CF488@R_^4O(aC<7LBM]R6-P90VN\Gg9
,9S/&^/^A04@[Q@R[WMAUfeb7.+?O9b>cI,8GO?Zg^P4S1A2<1).Y<XOOX2dV9eb
F)3?L^-9MI2?0M;G8PC7H8;YV1_R<MTU:1:_;bXU5I1NIFVd[2=Z)dAAANY0491W
]+dDc<LQdWg16RAOP?:\54c@Q,E>_.UA^b/8TPd/54AQfR>&<CgW)gY+@D.2?VXZ
_-+T&@fe\4W90A8O_B^2U/(T]Gg?45@<BTSRdJ/:2WT8R+HB_4-;PbHS,X5;2KR6
(G2529-K:f8&.W5[4^^:g,V6H1^<<4HN/&XGEN9DBdC?D=aVIdcO7FKa)YLI&JJ0
#C+<Pf,W/M,L1SeaUa[TC[YG>4H?&J,\<-Y,XM&HA426eJ(3A6;aU4,Y.4;<&cYE
+3#\?)-C?/;?19V0D6]4fWF:E;bLPfLSf^4/+a>7Z07OBI]2C-_#Md<WK8)>(:Ba
-.XNf@N(][e\6AY=F5H<),FLH-4]11(GS#1KIaLA&BZ9d4&BTJ]/HOUBf-J-M-6[
JV59UL9b9/YQG;I+.PX_13RVA#KM\^<D?>38WFb1_+/L^75-59cbG<4?(Afe.;A5
?8:(X-\><\Ig6I8/C9c]U@QY:Q[g2b2P?;,0_E^Q(3^):2)X<ON+WVR7P0@W:<b]
bO[f458QL)S(,MaR)3a.Z#c8cV<[Ra5JW>><.QLB1/]\Da#DbEQ3QG1@1d,R6M-[
>PfXH#fAWX7-##OIAUMCKZcGS\V:D@C)&L:]A;QLU,P8;<eH4QS?dY)N/=A;R\Ba
NC#d,/NNSP[5AE[bOWQ@>+CN5g4)()V+_1O3WK?H5<J_,VbZ@HV9,W;cR?W]fc60
T(>VNAZORVF6?HP=7EHV;9e]X9Cda<ReRCL=#1)gN\V0Cg2WHd1M1+X0UeXHB=U0
b/VUI+DG>?91e:[KIHSV,?1c_DSZ<68ZeXgO(E)_f>57_9(50,@RdT7Z0eBTINOM
DWc:U4STVW^@[fbRWGO(c/O6O^(8adN_,HbDQ@E^6_OEPKTW)CJ])f6e^K8SPdc1
M,J9X=+R@f2Bb45,(N.N7,Sc&GY,eC@Ze<&<:_)[gb5ZEEg;c0.?D:+MQ3=>QD@X
1DDP8.P\\7()RDdIaCdKEc[^(8g@YPG,=GFg[M<>g1UNWY:<F6C4BYKKefEg.&2<
B3S#8JDBRdY+,82J:9H3G9@Ob1eF4I[VE=<W?c]FU^b7P&5bYcL-#E]BI/,K#DEf
[,_DMDa>3RKBZ+d&@c^\BN&)H5@dJXfc/CLg,dJYV764JYNI._NC\,a_=5RZIT.?
Y,5U:;W+5\DfC6b(9?c1e9<2,7(H1g+@R5GSS]+c-P_R.X/;dMdfGSab.Q.S)&\5
YdZZ=aDGa4G/dTg5CEBARO78#SO\J]2116a_H]@[cZcU&F6+/Yc@9C2R?PHK1bRf
SIU<0I(=BA>f_]T9[D_+OM_5.9bU-N2;5/3FJC(T1:QH9.&]@e)-ZTgeNJ6+)c,0
_)aJ(.)TKg1D@FMg/OIZ.d1>,+MK(7B.4HFg^KM--+Zdd6+J/YV4d:[Zd:,;V3)G
O4WXDGJ_<A5/@f\=>U>,=-KO[@CZS(:J6IOFEZ3?B,]OPb7T7+P>M[(B=3?/I2+E
#BXa^283f<COg1_M9Nd>AD8/67]L(L5X]V8L8P7Q,+LA.ScSXWLN8=>7JUObPafb
QW-&9GJH>C,L@WEL\].fH<GX59W<>BV5[(Y&F]#3AHb)G4,[;;9)gP05?[gZG6Tc
W@(:W[.?I4PGL,/fXf8a#BR#:@,^@.eIGe84dN,2Q^?CEQGCUS=c(H3#8SUf-#;N
9#,&;]#TBC6LNW^8<3:[)E,U<a>Ef[[e.]H(02E<>.3ec0a]Q=Q]ZgT@.T[bUCAe
F?:05=1S7HSCW(KMg9G_P@(=L/XcIR3=F8_AGD&F-UGMScB,CK70;)F2/DAU1Faf
:N_&?1NG80,PIU-S<4SJc[=.GeAPUGeI:5@df;QDM<]BM=D7VK.YdF?UQN3@M,WN
1;O8(c;9LPG@\e]?T[C#5DWH(_8U1eY8#-&WBY/;E=?W01?Hc3H02<LOe@Ag1a0R
Cg]V<ggEOJ&HZe[<ROVW#-FL3T]>P8IYR.OI_?:FPY6PB]L/B=8df>[da_]MI?;2
3J38O(b1@N3I&IVXH27NVMf9;2XWcK([<G35V\NbX_<6&Q_T?;D;3gAFV&(>Y)&d
&T)#f#?MD@;W#S:N1(:)0J-VF3OFECG2/gb9@8<;-Q<S08=Pb<gISUD]\C2e;4>=
Cf+5b&RFYM\a<<6#8M#@GY6R:&:.V^P^Y^cVCY)F2ggJ\YC)9Xe?6V#.WLbNV_Sb
g<5U++A@>B@;#47<Fe3RIfe]/MAf@F,5Y\X]59b[0UY7I>.gb[;Vb@Q@S)9OP39J
L5.[/Oa>D,)D9@f2@[W/TH3UC+PHUX:+;+W[-&4Igf&XBfWP48GT1eS0LG[J-G.>
#A(..4=XX[Ug&@S)OCgIL?M:X8I_Id@<0JEU7][R^Z_H:IT=283c[c9V@AIg9F0X
).^\/RQL78LS-IDU)?3-V1]-1_D\#b#dSV]S&\Z]5>HN\[R;RU6TW7T?;74X_C>V
_Pd8DQULNe+A9Q.#XOGHKd[;-W8)aBVL(LZ:E7V+8eB9;d36][c[G(C6Ze>(@P>N
Ha0X&R48C0a\-C+0LF:<^V#-g,C+JgI:O78eDB:CL77NLdLQL-UM24249cI37fHg
#T-c8EDCJfCKO.\BX]_d7O[Ee7-&GF80&+eF#BT4J&J30X9b4X7QR5=L]=L-]3ba
\VN3&Z01J(>Z@;BdD\fC.Bec2J,,OZLG>=/^DcF;X9f3DR=Z;,Y(X8+c85SSNN4?
:OX1Bd4O:eG<)CcN03b,3E3QUNC1;-L32DU:=g)V3<g_/_?d(D3+98fbY]9YYO1[
&#5db\WSLF,c]KaaDCceT_-8#FCbF::3MD4KN,.&fO\7gWN:,^.:&2\]9Rbc\FT[
.M4CMVWS:efO0J_bPcZbX:gKeT+PRf\?B6FRVBPZ03BRP2gCEbLcc,e^[-M3^GNN
1KK3BX;Q88CdbHBNJ]ZE85&Wc@?@KYEJe3.&SD<E5d8/^0I4MVGacHC:eVLd-LF/
(;a8_D5KBW63F5E?_PfKM,A@gg83PPYYZ6#S9cV?E\J,.FPLP>SZKN4=[QW_TNbQ
gQGe6b_HP\I7C^;g?[4?7&W7MW=,2O??-E];Ja&(0W7II:EF,VS:P;ML/[[QL59E
2\DXBSG:4<C8g[HagF8PB:,GFcQ<3N;(_-b?.C2eWH]#LL@B<NRd0f.>.Z&gU4Wc
M+;_,^:b-b+@>N?,dZK1.R=[[(=/]X[]bA<LNf@6PVE#W>CYCVaH/^SaN=F+_\V:
1BV-]MGP+8gaDM4XF9>J4GPW\PLdcQO,P2E;Jd1>.(:=,L^<5_ag,8g<4/TT+e@0
eQf]_Z:_)?WHU4^5QLRN9g_>O0Y]?a6N4/,RB.8M<ABdCTXY_\NISWV9I7c8\:L>
RgH#HF>gd.#&KdUH[+LPOI,c]gMRdYgB3Z]HcTVDGd>LT#9R?_9?K9UEZOS4K<G\
O&FT0HA8;f,MbC<9+06Xa_AC<?0Wc.02647/JfAM)MMcZ?E5B64JHR>JLQ).6LI(
gMRCWa=RYR/e/F#WH@JN62L#d)(K9fK(QM6(U,3gPeXW\K<D(<59YV8NU684(gU@
.4&W^S:[HRYaP?Ba@d@RR,^=8)@G:RH=+YY^TNL_M<La)>>[[@=4/ePLETc_IF8W
U/B1#e&\8M4RUgZ5E]5^I4Ng8[WNd,W9\GZMY(_J,SS?[PbSYK9@3#P9ecY-4\91
LC_:(89E8YD)?OJIE#H3^;RbA<f(+EL-bO(Hdfa</M6EFdbf>8/8?AM>&@^_H[a0
^[-[(RL4G-KRZQBXG&3\B]HB3D,]GPM,P@aWW\\6KR,CIc9U3OO)I;UVaVE1)(aS
?K<2]N9#N]Ke@,]82B-\L4)0MLg<PV0U50H=25J\]7c)T0QHJaOG9Vd,_Ye_EK2]
LgP0g4?XfEGH&gQ^CNC+e/RGQ3=ZH_UBGIQ.^[Z(6EQ,f=N:&^FYLfS14\MYYZO[
2gJ]&#@#4B^QQLZ2_X<?CQEQA_M2TP@J=,?WW(=[4^;YEP)0-YRZg;)NdO\VN:.#
R6R#K]f:BT=-_.ef3Ga^WTJfMQ[ZHga6&;UU[.V<O_7X97R/:/T=4e1.YcQaK[SM
MJ#Sa-A3&7]G9BT<bRc39F;]5/aG2Tfb)dHZ=eS/,FE)_CD/c5YLdHR_(S+D#:P[
a3,,0B\74=FI=,P>QN2.)H30CQ1)-?e[;gAZZ3\<Y7R,FVHAe(eFUSD1.>O<ARYI
[TTFJVB>TddXS]bBgO<[[SeEM:IX4Oc&5aEcBFC,SWFXA=Cf0AI<6Z)&.3CgY1g:
Y79_].V+S4#+?6CK,=U<_\AMTAR#cAXM3;,X/=-GD1&,CZQ>,b(Y&IA>LPLQ/Gba
R)bfI=:(9:Z#--V/dA^34NK0cSX[f)&T:C7fb_\f8\IaWX</DDRW/9A&HdYT&Bd(
Z?S2,O)F\Mab_62<?7+;KO#fLO@<I+[XR305gSE1EEB-B+a4SaUe5Q@?UUJSc#TV
/dL;RRCX/K&<,;E&_FXD;cb).8E->QN\B7IJfMOb?I74A__<R@,?IW&(=2NPb82J
aMO^S0KP:)XfKQ.I7b69YN;[[<K8I/X+cE);Z7VSNB0@ba#ZGJ.LVO+g^BRSEdE?
6D)RO_\9=2Lb:@<PY,09Y[-8ET&4/B_8_f>X8e2fHB)fZGH(ee>FZ<BHOMd4e&&T
T)f[VS43b385DMNPRd@KYASd3@1HA@1ZT/]:EZ57)f3R[Y>YcLW>@Lg,aIYT2@F\
9HA>KP])0K>#]PEN,1)<&=Z;aWCU4:\:8>3(@e;S+>9gaBe9:HW#4&,Z7IUS2\5_
+?;W<^a8Ae@>Ug.1&@]G6;(O=7@^W&14J0P1S1<T13<9=g@,+009(QKWVa6Nd^d_
F\45f0[c;\/Wc[+9Nd_K>2OIN9BGb])K>JU9/+P:D)-L)L&/L8;SNRDF46ZcW+)B
SHCMRNSQf7A/c(=@]O@2@B<(@Z)Q5&[1:+F3fYB7:,DWAG>4+J5O?b/3225_<XN6
;>]E?@Y;A,+/#\9Ie.2,(3)C[P>PJ<gVfYWBD-VUW[CJO<-3@^6E1;7g?H5a&3d_
U91<VSg.bg&IP@+5W1O5aFa2f.&;H=>N@4;ENY&b/.3.U+_;5/U=2D,Tb]\^FB<D
a?IZ1N_@e.P14Q9]@3>WBce3#F6S&DM9AK;-K1JN2?3]9<a[T1&]PGFT7RRH[.>+
LeTGAF\;_PFMZGc_@+29O)3>>ge_P,K^W>L>D#3WM3^=WG[b2(:)?BE<]WQ97Pbd
0a>b1H:OX=+NO\XV6XI+D,0JHHXBSL8(cA-DZR21b3LK_4)&B;.&?&-^[e#]=<;S
&MZ4.+9-SMB6g=21VecW=a&,-Y^;/>QSe&\?8O\/L_H9(FaA_W1[_B[Y(MSLK,&7
A6EH@L2#[_VOFS;5:7F8YEFFF-C?W?RG[H],&Zgb0FV3Zg,AD;FAAbPYNH,:[N^D
G5N0S;7gO,<^KX,5\)LZ/F\9&BO+AgT=7J1&A#Y-1R/FcA=@>.E07J^dL9=>;acS
3)-144JV_.^OO)c\0X_U7-N@RT/N0YC,=Cg;eK7&6]J\)O]_1-+IIRXT+T)QUb1P
OE38.,+-;\cC(^:_-Pf-g131+bfJ:1M,(E8e(S5&#dg/d715ZG0EJEGKSI=[T/XK
DX^RJD1EG5WTE<c>_e;D#W.YK3)YM;MDYf7#<Y+JBZ>2+]gNZc^@]\LRB?G)+XRQ
]]DN:]OB5@?2O4]1G#F..B_;;+<Wf8?:DJRMCY:aT=1^X?4)G.P-X_>>ccf/F0LV
VZT?=R\;0S-c+dUZTeb)\#5,IfZ7H,M;D[g7)8A=g?0B-JgTGgDb.#cVf2(V:fR]
-TEQVG5I/V(NQ6Q:^E(ACT60aTS=:TY79(\WHaMP+URLCZGaWC3++-75DNB<NBT]
)DT(fgNL_4BA^b,-L;YND<OUQ^(TR\g4g>GX/VD0S2?H=^.0cg:OI<H4e7_OH?aT
->Y(?b.Rb+ZD.8D\B0e22TSg-6g_2+;NFD)Q6<EVUWPK[1/32(4+dJEIADQb];3S
?eXT&Q9G1\c-9.;0T96)04bPTN:fA[8,VRX1NdW+=;FgPRE;G=2T,/&_V4S[)SFS
6/FEL6/TFG<G9P4UFUe]WGc(\@I@^L(g:a^O6\C-Uc?>UKeW9R-B.^=(MZ.VSfEO
(0eGK)V^=;7BAX^#JC2d;L&A?Y6GH+#M-E5g]IU-X.Y75-S)9I)BJPTEQ+2^fJNO
]MTC_8=PY&C]@55;?&C5PF?<D]VbQ4EHU=E&[\6cJ\]7)76dW@3Q.Jb8GeN,#0WX
/]4dM+<>D8W-U/KUK\CWc65(JM.U9c6-Z.,2Yc;aT6DRCX+8S1-LDSU5@cWK1T7c
a#1c:,dG(d2WaRZSf6\c1+Z7<M^]QE_,Qc1gYeDD.K2YTPS),aM.&b.c:Gc/=eF-
:V1ReB+,+g,e/>c4\HMM&;f1dg?-/KBe)M9A)ZCR7^_YYX>[7F7U6eIHIKfdUU>7
Ec0Ce(Q</Z1e0S8eCVcN3?E=(c,9C38gf@.Q\++f=4B/RSB5W((acXUJ)0F_+//?
:F]:9K=QbXRS^?Z]HZVPQ,Lb,ICfK6)5Ga)R,O;\W+D(Na(S^H\UAL7-/X6NP:_\
ODH]6g044ONOI;1LbM(QR[I##\Y>T\[GW>^K9=<A,>SRQWI,Q(O_GO+X&fEXOfS2
]EC:T2W^c]EYfT5[BQQ/@e&D-Gd&Y1W5H[SM]ZfP[(QH-<WeV.STP7UB=(NS==I6
@-\])Q:1fLTFfKc42Qb+=@PGO/5dG55T3ZK7agR(,gc[@:6X8AYC+9XN?T[3f0NC
8D&J:AM;@La\42RWPIb0E32bLLB_ZGT9=IWU.ZL-GNOSJ.YR/CJ&1)ADYVfR,HH0
@<GEMX]40G@/TS);d_CA5K^aVc2Y=;09^#bb)SJ+&=HcR/+P@1G4WQHT,M[JYHTZ
[(S2b0:FaRL?7_+7DLL5d?.U.F7fFEVQ#:<3<ON,8B6d<5PcYF+O>\MUG#_c:eL5
16[:d-gPM]R2b,e+P0=B6#TL22VV50DN\[XSO]A]4RYXPF?C.8EI74GD1]VJL^,]
\X53Wb4OC8JQ35]+[(RM/e/G@+^9T&-89C,e6>KA#_+\&<&J,.)WC76G@G5TJddR
FG9MQf.b/W0QODc@67\83_M9bZ9HR.+(PV,6b2C041@;feS5&B?Wf)6YYF^-UEg)
4ZbYD4VDO&)Qd=4c\H??gMFVKIITSf/CgW,d^e(,X/eB<+=V57IZFH5:(T<-;(12
(:3Rc^WLPEP^&ZXGEPI4QLI)ES9HPVTDdZ>TP)B+?eEKVcf(PZ>cL\cIZCN[=J+g
;O,K6.G7L+6L5VR^g=.9RHB]G/23-N3=D.0Z4U<B1a]>3Qe,(R91bOBT>SQVHVfA
J1A^;8,4Fe(b)e6?DX1F7],LgAGOgV[Z</06/g6ccdG?IZ_C&eL^_8GDOb[2AL75
aR,>[<[@\^5LE:[T#U-:d&:<H\A1E3:a.>APJB9dS0+IZbO_Q9JcdVSAZ2:@R60g
SWf>[g>+>B^92+E_LQA@_<#]QdMUZ7b].C4QVe?gI;DNAD>7_e#B@UYa+6-,&S#c
<I@7WND,5,MeJCR0KGdPPd0>A2.HFPJ2.V^.UYL2Ka_bLa^X3RO1D1fMY,NNPQG1
X+7eUNKg>/KS#dY1H9?K3cP@>HAWgXD\H(=c<(]a.g[XAaEZH9OV#N?&I[7XR?=.
.1(/AF/T\:^91&2(WU&XA]EUN_2dSZX0ZCC(a]#:H9BU8aTg@dP@]O9bcd26-J1)
T#@6fD_g+7GH]aOULV,OYLRIc:HbQTfZY;2O/LDARO:8SXU:R3fK8.LO9AY4^6OF
_O6,(\BEY#,5Z#d-]]>VfM5GA1QbU9Z7/cNRZ2>eA7a?V7DS,1-PcY?\[@O-CX;M
16(3<4QWQYV9;+F<a]NgNd/FH:RR0KIE,HdC&7-T7H\(d&J?A_OMbbZ@46Zf(8K7
5\&b0+?T))Webb8N//]Q,DM-Z+OW3OJdS#<?Ygg@ZFIAUNOG6K2^_aNWL[O?L-91
UQURR(1X9(5U62\+U+N<[W6b0J:]XG1YgJD/DR7D5+P<DFOR;>57MdKL>Se/BXMH
PAE8.M2L)CL^RJ9Ib1c]\6/[)e(K&[8VSIUQO:P/.cEGW4OML=&C33D?M-HJJd84
bZGEX-d8O64-W4.LD&NZ^<NS1PVXY.,)_EVM4._UaOD0=]AW^KQ>4OGFPI(9C3M&
Q;KF8LI6f,774M#[FWcTeZ8eBD<OL=^#_#[VKX;Z&&6J,L(RT8):9=&gS?.;58E+
<)aX(N\U>XJef9CD.(8^45P(+D0/I,YaRM(#LQQ9^P6gN#]CL?>,dF7_B?_F+P#B
be,aK.;>E[G4;:J2;+,7HA?X4L[?7MT5U&XR]PAIg/-@DDg9I<Je)+[NbO8bAB]1
D=WV@_A^=1RV\\:-E/B&IPV7?NWNMCO4OSe##3TOE:T+QfB<K2>9WFJAU-IIP[J;
EI<43UT&I\18H#7W>I\N[H3TWP,^[0fdg]WT23U7I_7ff#<]X75@SEYCV9S_H).;
S?9IacQZ5-UcZfS-2Q.GHV#/FY/L;+c<b]<IE5Y#@<-g.)SX1\AfMI2JK?ORK>&?
[+7OE[UFbG5\3GHgP6Rf,]W/gD0fUW1ZE.U(0M0Ld/dX5.(KYb42bD02&9/T&[2M
Q]P9>#W845ON9VIXFK;L1g>bZe;U\K72E_g>Mf.1)TT5LDgBPJ4B?/8HW3XHE]))
):A@\3RE/F676D#Y9)(<2&?&6.B;++>FQWA2Qf=EH@7R3LL.J>bWVL-EB\RLMDZ,
/J0;Y/3+@CA\1F/=LE(CRP,;9faWOa_XDWNIGcB:EJFdcAXe.&Cb&YLB;@.P7f;f
_/?=M@AGK<JS.JB]@?52F?7f5DVSE(2,R_9#R7[?E3GCN)3J8\>dOd?\&]Q=V\[?
-6VA=U&5CO]<JT9<He5[57]UcfC]adA[1EUbB+4B@a7;NQ(.[2e>fSH0CG(?:eG;
;O@@Eecd=H+Sg96N2-]N=fT6HgWZ#W:[e9.E,V7Z/K;=O_aS9HQPLG4fR7##A0&=
^9RZTO/VM&9?8H2g4K8.?+CYZ5&G.1M8E=@H,7RRLJT07QIf9/396(9_7XB4&bO1
NIc(SZ9d&)@XBGZWS+X=:M8eK3d&dcVc8YT[SC=?YJ1@MB_]43/(R/H+Ub8)=aW0
<:OC6P@2OQ#^O_SU28Bfa_::-_5Y#>-0\T227WWIZP=<8X(P.[6fMg=KgRM\fV]c
N-\4[DHQ#_cb33?M;&7HdU&_0<UIZe4D=F,6[E7IaYe>WW7,V6XB+K+P.+HXJ<,Y
-=8b=Q>:SNb;^K/S>bb0?PG.77S/04EJ;b>.6^gPg1X79E7X^g6U]9Xb[9\_#;[K
61[cE\Q(]9[TcUOb/gd7Z\=9,QH1XFF2A9Q#:>IAfB/a7#[/\[eC38\@O]gNTVUL
g&)(5gA2/<_/7#5\J-&CTC)a4V]g2JQICOR>A4W5>PJCUIJd6A+^[7QB74_Pgb(@
BM#.4.0\.M:Re-7#IH2HM75K9K]G>?>3bReDMX05U49#\AMPMS:H-/+QS?,bJ99R
17G9#J=8>Y#\2<Z8QC-0\4[=Z@U2N\)6b@-)CO+@HKU[H[5c&b#186,cCJ3SJ39b
#Cd(L7#9J\;BIB;32?.&QJ4NVGP(;f?5TVN9)7gKGb_,;IJ:0+F7O3MW^1eRLLPR
cFdQb4=OecNMfA.5S+M2[7I9I[-a-OZ<L)EJ^GG-PN(W#&ATE4P0I>:(V:6eQ7bH
?+R8aC#,TT:73[Y4YS,^J\5)92+L>g+>QSJN@^KfdQI=PT85/MBKNYG:0V<#1)eH
ZVOQJGW0[W:[KJ2S37(71dc4^_LT0gXVHE792WMa7_ZV^GK(S@#T-8B=0bfU0ZLL
#II9MA;7WU:>VM1-dI5]>6fI[-XBQ\Y35I19O+^^9I\ZV7I]5]IK<[,5GSSOCcDf
gL4/dCHgHGEf7?^^Zf+Sb\9KA)H+4[^5dPdW;B_8L/45[dFQXCXcW>NO/2A3Q]ZD
QPVCg>M;eU@\/.a2)0P\O;4@5f,0EFZ#Fb2H190RHAT5N9=c=e_J)WC,aeSOeOKC
QbK7:OH7;7V3CRG]&;?cR\CT#J4=I:4M(=CNSNMW&2]>?=,a6LY&3C5GBUYOa,gY
a2-PZUQ93(7J=A_O\0S9+JB/>7QCcOHKeUCb^K_X5G^R>]c[13]5--e1#T6\R-42
GC7(dUQN::YVL.U^WQ=<>]Vc=AE2c.gV[ZCGP4]V[/)4B/P:X33AMVD&g691QP_.
-2MgAZUHM&P@]F2CGO_/F^84ONc/4U0@F^HT)=J/,V[H2>O1-T50IY:M,V1ZH(eW
Q@0DcBQFa^FJTf7Q/QB1Z7I36L-??BJe-A;UI[PDEEOeK-9:5DYYbK,d.HP+_M+;
G<L?#,@=#&gQ?^.;5=Ke=Sf>OOJXZ081@?c]GJHf=4M<3;5EKd+/@S([[R+#N&3#
L7VYA;_Ia2OEVX9-Y.1O3fbaPT\RXgE2)?B@3AJ#N[YO>]XA8Q@([4-5+VHg>_GE
MKCgP89g8GPLb7J>.--JbOUW;eAFGM)1PEQdYN8e.8[13V--INK3;ZPL\W.MX<S;
faQ#M<X_,IL1:0fX&>f2Ce#+b0W95Z_gGfSUUgPJ)49T-/b:V_M0],7f)/1=84S\
Pf3.e.T&IAFW4R@=YE4;S3ga\HcRG;[bU:94-K&b/:.I,Q2VAgTJ1E#3Tc@<H;2K
<.D]8L^Fb^@a-?]Rc_MD+UBXTf)ZeE]NQRS@V&?8\V=.XK-+60R\6,M3YQ7#(035
Q1VAYf3W01+KB(gc-4H7(+M0FTZLIRV9Pa\[W&9g3F4<8+5:]Y?AXWG]<=f3<TGL
:;H/30Fe^FB]d[Ygf_7<7EFR]U,<<F9:Ebb41#bATFfQH1H7:&BgXG(\bP61,I;L
;f9)ISdc1CG:Ue<YbGXAT)61a\@9<Pe1RO-5ZK4d7dMI(5>8V@fQ5ST>Gf<DX3FY
XC\6@^fW,H8C&B>-F69HZS&(c17EK@X7e[)7-5BH;C>+R(MGbOZO/dX7gYbVD;^S
-=g+<F=81YF;bEV]P(H=6IAMP#7\Y>]\<>M4HN3F6\VcFg<;-+bT63;g^^3WYf9^
2E=Na2&2V80P#@=&XB15ZBT_NO?0HS=X04eW)J(GFA6,f[F9Ib=_H[W,aT&XD:(c
@@^8IKfcSH0ObW:JY\P#+G^^KR?KFA.VCDZZCP2X9\5B^-\#H0I&ZgG9[:/0(N=8
CCX>\XbeD._?b8dF>CC63AJ\acBR1XN/8W-/BKD14dd0RDDZ]V,ERO][7A_Q?KJL
AFPS(]e18@,=4WPAR_+]03U1+QF\>((RK]HYgS[UTgYJRSKCgPZO5#6>bN+S8L;O
gJ:2B72963(X83<g^\&AT=OE2\:Y\X=gVW@#661?a/=P2]XU95UcXZ6fL1HU-03M
-<fEUKdWe;fPNW/CIXHD._9a0@.fQ/+FYHEA5K/GeYg^((9)/-Bg14Z^<IQQS5?,
V/]^((2d]B+YN_UUY==FD_732C3FXYCA+0TV2dZ?[DRSMZEf;ZT/X.?fSEg9S]3G
2WB8T6S<7.KAeU-T54@fF[9<D8(db=J/#ReO+4#IF^0-,CgScDfb6P6/0X]ASXaW
V&.]B1g_PcZ>0C;<Hb_bg6<2.HaaO/S30Q@7..@\L.@=>EPHe,QX6YedO=WaTTYB
UL0T?4C1X?1Cda_(dQML_DVW)\PR_1aa,65VE4+bL&1SbX9C2Mb3-H?-Xc<MQ.#J
=)ZM+ad]K01;:L(F]aUCf:KXV9Z]X8AB/2:6Y&b80A+Qa]Pd9MKLD3>.&PJ,<)ZG
NNOZR0>X[JfaL55dEc@4K&).I7gEO.a-\=_J+f_PQC)Z]P?@MPP2(#]NJ4MW:OXd
FK>eSX+(1E5S2YQX:5FIMQ1a3S]JB9\,EQ3Q16(A,6K[aY-W#WD)T&L^#f-B-&-W
SL\c_YT.:HA(U..F4d@6J#d/V2(<DKf9[.(NO_Qf8D;9WD\SeSHS0@,AbD-ZDE3]
(2>.@1e_A0LU)L0&.fF,5<D+gg;Y.BG.NJ+I&J;1-cd6W=(TVcf_cd)H1eOd/..)
+3[>BMG\/87Wg9f>g)1Zc3eLO#QF.O@\6V;EUF/:K&:PVH&O>P3AbGI0:.c&]P#7
5:d,RCB264VVdL<EVN\+;S:HOE4E)S-6IV?b3dIB+(0?/gQ^JFJ4a(NIAb^QYGO7
]F:QI@g\,_b0Q<<7W^:_?\QRd,cGf^N[D9\JK7UFL0M3Z^Z,;J3BKVT&5A4K,4;H
VG+F\WaEXeDSM]>\f<SLH0\7B28^V2Q+D<=,DRJ@2DI)5Kb>2g,gWgROZ9#+M4,b
gCW-.1ADS\_?<FUHE\;@I>5XF?IIbFcQJPQW8>V[89b:e<);\U2&DS=,GIII2d8[
?g:-[@ZM:PA^9K?Y)K5Z.XSNC/aG[>f.>G?251YH>O/9f:59a,5cS;;]?K>@Va?2
CH[gT_,Tg-WB(F/gHXJ074?aQ.54[4CdBPJCW)b\@a?P,3CONaGa[2fG\GR>ALR9
\&dH4KQ/NJW]a/H\6,gf(G34-HFC&4cT+M[1+dT01\]9NB>G+FJ2;bdDEU]P]4aU
JUIFU?3PXaOD:DW?&Z]R42<G8U0.8>HFU)LPO=:<NYO[J.G+b0R-dG092SX+,B2]
R5XcP\QC)7RL@(+#M]I@&-3[=9BgK#dHKQ;LF?1@&f3):6c3B?A>dg[WaHU-#d8S
DOUaIH^Y/X8af<4I1)DMTD(F5R8=F&Y#COZAAS@=M]X#(3[,)K3Tg4-dM:-QER(b
(E4fb0ABdgYg9d<&@O4/0T=_C+C2Z;;aY^f&?c\>+GT_\aJZ8F3+GcIQ6^c?Y_/\
&83PbSD,Z7MSf>K05WI@X]O5<?DJSWf7:GOOcMV-B5CA?<49\N(]&a3:7FW4-7#a
<1K,2a[Z@Ee,_U_:-2b[P6NEDCPXUZ:0<7?URF?R9AMc=C4^]WSNSf\MV]Vg-8.V
\VYXF.ZULF<_;3;<<O).;gJ?CXZ;?>a(_e_c7(IPSRZf3a],J<-5c^#K\D,W;La-
J/R4(-KTRW?V](^1f@WdgT#RC2#TH?+91Q,@R9CKG(SE4?I<V(1G(@O-d8PTA.0+
c&5F7NG4WAbRF5Q\-X25YY3gUXARbL-26.L</b\RNb+6H\>&^2GJV:;EdY=SM<:2
\,=E2Gf<T-@WTcaDPP>ba4TDg#RCgWTA>(Ea?#Z>\>7UM?)g@J\/:D3#4gdYb=\N
H:E=C_US^9IXEO6F&4bB7[^/aPaV:_ZY3B/_K@5>871_WR/LTGC<T):;N=UdIgJ&
WQ5O7#FGG?@-3,G&P?IBReI]CPEeTVO]<HZVI?P2\ZY7OS7E9H23MZf]=KGOKR-Y
3DXfbd2.M6I\QF.(U,:X<E3->g-.:U_[VBK;/<@03E&>KH31]B6DeOEX#RT_W7g9
X]M4VU:M1F4G62BKVQU2-XB=FB:;cTBGW[eeB4Md;,#H]\f?Xee+&8=2WY.WJU[&
(XB]ZB,bDbZ(,[.KQE;:A;7J.EdCL&IeAMZPVN)0P-0Z;ZTNAbQOZQ;>)faf;1Jg
/_D\4=Hff:M1_P>IZ0+0./?EP,[^/,.C.<-+BeMFg@RQT/g1EDbI++KIKM9#dBHf
TY,S[DBRO]N1LeTd_DP#fR3Q:4,E9bMcJ9^E-f7\OQ0_853A,:7YD5[FK9#(0/gX
]XC76Z/X\KeH4=6JY5VfU^,Ue]G;T>H0RP>6]Z&7YT4g>S(TZEQDcU\dDSZc#f_a
-=PV+U6OFD;W9(M&<C^<[E61-NBcLRL3B#F7PO4.]/+QN\3E5S5@SN=&ZJLQ@?^;
?ebLS^+.0[I?.&7MEV\)1&QWN^_4G0JDRD#c<5/DRT)g:<e[&&RP]W;I9/g+F_P(
Xd_8&R@<gg(E[)C[3QJ^f-VTd,e4Q)U6\F&B,dI),#_&^ZGHf=++#5(U?ObCOHWd
HNQ@[-TJ#J4X3:e^>Bc11d5F?;.g@G?_Dd5Kb>6JNA->H@)).#(]_?Y(GA0O0R4]
Gg@gGMD][+bD<VH3a85&D,E_NdB7VHM#ZcJ^LV/G079M&LI564.#^JeKVNFQ-HYP
G/EN<U)WTI=;&2@T.OB<PTE4W[(&.?eV2.[KY3Ae?#IRY9>51(+Ya(B5CQ)Y;[Q7
+SXH79^?dNHR)REdKD5e3AIQ\LgcTQ+Q0VT173;eZX?McM4_=9+D:6?TJ#FSZ/F6
=J8\^XFKGF@<MYeK?;;N#MagEfTRXWD1A&MdJ#X&M[R?a4.+:U\NG(,S\B>ZZP<X
YG9g<-V;gG?.<NL]S\6.QPO>:.GLXAd<LY7635f:I-f>1PQ3V=CE/:WOQG&be&<A
P82gS-&.JCAM(@^Ga;+?7VBY7L+c-a^c(E\EJ22dO1X@,&Cc.3<@YTSd6.#M#Z[:
R93?]c^JTc\L\0FQDC:ZB10;;,7RDY5@;Q+S/M23]Ce^cBUcb<Sg^../;3]9OFSJ
1VfBfVY;eTH>Ga<Q2#C4291&#dQ5])LUa@0P81GgMP387@RWQ-GVVQPaKUeRaV:L
bYN\GR,9OaAbC]0<<(]UL[e>#;D-6eNS9QeLCfL]FZ?TX,5^LGCZJ(gEV^DU5cWA
&;Y^.UQ40ODK65N_b66U1Y>1HB<&S(8.;Y.&-SP12HdgU4]:/<[Kg=ZK.^:UJTd2
VS,a&E5IVLd52T7719gBf=+?J];J<f,I1PZKdFLIGd@e1I7dWQPgNY3cIK66c(9.
NCU1]K?aDUZMC?B&fT@G.AC<E]DH=-YV4M7Kc#>B4N=2^O:;65[/KbRQ=B6I1QJ^
JYe:<M+eM^>PW),[=@>(CKLJ>]E=I<:3F?IePCd\f8.7g]V@^/G\CN5UA^^ZcRbI
<U^WcZUT5-SBJ8(e34SWO0\Rg/RM&YYB&P-9/1C5+[X_d]O#83+eANT\8gEN1SC-
J8C7-9e:\QBLGX)g_D29Ke<OJ^<:7&,\<G]\0^8+13X]KYbYP6877b04S&5a655:
VSdTD.HMD_:8+TT8e^S?W>396LbdYd=9__FUG&E-3gaASIE\G+,>@E??/b^I_f.8
NJ2\708J4_-2[4..c+^WLCGVAS([DZ-HZ1JK<,2SDML8/\613AK@+^KB2f[f&9:3
BbPJ,\VL.:H(=2MQAU</.cE78bLO[8M4Q#O@BR-BTHN:d)1M_Z2H9IM048X@4+aZ
);8Q^WV0V:4@OBXMB-<IH?c9:S2E<3<-EOVRH4\+[cXK&2,O85]E.OC(RH99/+YE
-.(JJI<+AdE8#(EQS>2+g9g[.2E;54W3>?_d=;]2XRT)W::\JG7(g])&O;a80HP)
8&>4\gV5Y.\_bE.9\ggOM<eH(6/QZ0/?/c)Q6QOHXLfCA)dg5^3aJ<TDBD34(R7A
SIb)D01CT9@db>),]:,:]MRR,,XbgDS]9.8SSFb?S@Y.=C<\I\TcLY-YHA3:VeK.
4S:Qe@(c&@V<WeT]=N^QDR=KBDPN]KUECP6d[/W,FP?2Ca+H+AK0@=7fK:+M0.E]
ASP0>HGOA4?UP)YDQ@8\06H>f3U#c&>B6)40SKA1?,<8+F]aL_cCHa#T_3WUEMcZ
+NJ:9+[d046gd]MP]fG0Ze)c^aU(Z-.b.YJI=\AR0.[#VC\@V<KUgJQb>YS,#LS&
RA2<8V(b,Re@PTc_Dd:RC>0XGO#@g(P]_Z_1+a,#MY6/V>OTNAMK;#>L]T/0O[Y,
+Q8TX3&[8EPc(75^ICa7+TJHW&@(PTXG.HQ1L;UT7aCHPE4]3JV]P<<G4\97T9d:
Ae9F?45AI#9QJFdf[L-T@PJD@CY5K5HeF0.#EB8@(5<5cY?@KEB#1&3;G49bcJg#
NC;d<5.&WSB3[058>ce\.Yd[@df@<e(8UZ@b@b/f,>KZ9J/S:7EaM/S)T_4\NKNO
^Ia^TaS@=6?Z7,;EX5FLZ#eY&.Wc[?,JKeA4.76>SbS--[QO37@R,@FM0E,+CKR&
L^IN9H]L[<@:V/bf+f\de6)Y4(8B9<1fe,R;5+DX_DcfB&g)X7+D\dZUL9cTfQ-+
[+DdO+-HZff6Z:<=55aH\@WebaK5I<@g4OD\Qd.01cPAH8+C36Z2SXeQ\b&Wg+E<
R0(b83Z+K-F1agXc2WR]Od)bU=43cWb7)e3YgAL954HV<IKU\Kc:1GEBGX]SQQ(8
BVTHg[JQ?O<P;CQeRZU_A+8@bXLIA>,d\^D/=0I-4aQfeF0bJT;[9dJJI+5F_JS?
2WAK8H]9:U_e(H;BK#Jb3=LZFJc53L,6^].e],_O8\A:+NP#4#Q9:+)W9)60)AT9
.)WcRY2\-_7OI5TSNFRA@O<C(LXLXOT8d?IME(gYAY^7g_L1A3-a;3684?_30#MN
@ZH7VMG:ONg,#PbV,W?C+89T_?0=&]K1+HN;G+VCB>3+G8&EYZ_FR#:X@^PDc+6F
@L1O7I5^#PDK_T<63>PF[8TB7K#,\>LR6:9C?)1BE#27:C5?B+6XaHIMG\O2Xb35
[cX,#0_TXPVB#U5@]R.U.VdYNfD9RN@^D:Y<\UGB\+73c3T25<V[1[2dY312JX=&
71;[H\^9HG_.-7f]E_WUQ/1(2,9[.DP&;^5Gb^fVA&)6-MEI3=P.3.<G.f\GB4[0
Ig=F(6J^W#R7=B2586P<U@29N)HNAX\6F,N5L7X8LfX5-7.VO5gP4WZ1TJ3b7E_f
TK4NP:=9+Rdga(@dEa=_E&=+eP1+L]4<\_V_@8Qd35LS<OaJcR87Ia1R=X-.e.A8
Vde^Z^E>C^)7/70O_J5#2fVY.B)K_A57Y]U7#S(KG#b<4\6P24b/:CE:4+MBPeg-
7E33];QK^#KV\C+0JUUe-[;2BO4S5GV/I1X5d+g?(D-.b+:M0.0?SaE/.5:f]\>L
FG[V^2N?ZfP8U4G+B5cE^JOgSN6R\#b-=:E+HTW97?FSX6Q)J1-1EVF+=.K3F>3X
QLRT@8)WRBFACE@3V?_5NK;f71NSS]4EO+H>Oc&NOH6^2?P)>P+_39e]AEHW.\]#
ZL8)dZgZ3148I2UUc8&0+#0b0R85a:LcL/.L?<9/&1\CbFg[6&S?+?L6KQ,SbOG-
^9#/W)Q8gV6?GX6.7fAHB.O6BS[G+&>OH0.8XZL=c39<bI9MX>F4Ea#NAQ]BNIbg
U1_#=ffVHKd_@V;a^3TABRL,7Ng7,NWH-0OEA\X2?A7FN+8M[IBR-9?=)2cL(MCb
[S5,A6P],+5?H/_,UF/g;G<aLM@B96AUB>:[@J05HC;M[dJ.;=g5JDXXL&?b&b#:
W6AR610+A(.aDPQ0L]Y5SJ:X+DVKKFCVM8BHC7598GUfB@2I&ES4+VZ9Ke?fW\)-
baN@b:1NVfAg\7<5e2C)+&ZMTY,T1<L,#J7/f0e2>DK/=7[+03(+F_(_+1EFX9;?
gC/UKYe?ZOWPGPJIf1bM.7A/R.Q7&[)ZNgANGccdF#1V^,_[+cM^/0(&2D0W^6:)
KCU^T2UK.@J<-2SeMC@8UHM9.5_c?LbOb_)C0UML0W8;4fN7/KgLSE7[ZeTg^E>J
N3W)K&NO-.]9,GVRfCQ(aXQ[[C-103/&0WB@<#,E&3EPGb(1M^Pf^8=EQYOHf?b3
F.XIYAW+68Q&//=NJ;@-=]GI])Je,d.cB#B.P@DAST,Ja1MO#PJ0d_fUCEfdVG,Q
Af,9NeXH3(_1gc;eV#HOC;\VV[RP:6VXeI^,/aLM903/4P<\(],K5d=>3C;_0U,I
:)8QM\FZ#XQ,2]=(:LC.+X;/1b#g<9Ue-HP+fL.fM&V3-&adPEQ.dK,<TDENaD.1
5@DI\dZJ/F7;R0P<bOV51WPQ=b+E131KeOF+BBgB:.N3f;\fK6b#GcdSMC_&4;PN
e^bI<QLQQO2Y+@Z.Vb>/QYUedRRMRW6(Q;bL.4I0[-e<bW.;fIR^g)PKQ1SP<929
XH]2C)RU>9<8[0FS33PXV/<4S8A)TUC8DXMcXJ<6F+4?.+--^Y2<30QP>8#,GaR+
GdT-@^(9EV<ZA&[9<,=;\E6X<;/N>H)eb,\If66),_D3>UMB.d)ga?Z+^9KH<I+V
EU1)WR(3V;+eR)1=c+WP:NQ.XLI::a,#K@2-?g(,W2HBBG^U+1c_ROF;J:@bUdIF
2HRWH+,AOI_W1FGU920d-.,;WZTMP(1g3]-f0(3cf(2(:,7Z\CK)PFIK:F\DAN&/
GMKbFc8:AB,P<8T-c]4UZ6;MDF^&08[IT,K1/b6d].Af=-/9g87FdS1).CGc_cF+
VTM##8M9d#PU460bee#Fg9G^ZRQ_F\X1C8>21[[>ZC\DD4PWGe6>b3]c=KVHdQ8@
-Fd28W6d0NWZI@D-F78(EgF@g2ZN<V,\=1LbS;[7&HQR7GMggF.4W9&dNa2U@9^V
997T?^1Ma8.QKYZ)A6AOHA.X@a+G^3NAL1W7X[^W^ZMV54V=96e=3TAca66Z&R;2
0=M5fFDUKe7fga5/gZM)[=T_&^648\QS7Ee92Y5<-aJ8RM2,6&[5W>L\If?3362f
=@X5Q4J]L4bOI-=<J[1?g\<DE0G(M1_7D7=e>5BBW2Q\9L/X@ddQ4]KC^d5.:0a3
)B;cX<IT-Y;H-JQ^2A[Q?E;YUN>74@4#&32O<d;P@+PI,3Ef(^RV@>9ZaB4+;>OO
/.G)?A1]4ea@KEBUH.WNQTcBbHcLNF>PEBI:N2UdV#e[@#YT;L7P4Z)Y_W>@@K.Y
2:)/>P=#&:P0EQT._,D/=7^H&/_,XE=3&-B36_>BfKFQ2_gQFJ6<5e2&D_b4.6VS
fJfCM;)WQ,+5KPR\E6Q&Z\^:ND7P=PN.+8R9<Z=<_>[P[Ma,84<PWS1L7cV&T&\1
JXM1HH_T:+dWEa/&^TC3/65Je9eI3RXT+g4YbC(]LWY0dVV#f>,7##,O#G2D-,0(
D4ag,UdgN5X.(4&07=g(#AI>\7E0-2ZIX/M@IUQBV+?>)Qg/=Vc8NS[bZE7:9W7S
Rg)Nb4B36+#DB\=@45@g?78C0LOY@P1#XR1\d<?<567AV&U@U1g3FcM691Td>e>g
4@W[BRKI.Y&(W;f_4O8#NO2O.;6R>TPI8e^<5BO@A=0W1\DdVIWgEWPKPU/VYZ,[
-+@:QX^THATeV<KIS\496&4]THSS&:ERIH;\R6+Q6II2+N??0YIQeNd?EF6+@6&0
)EJ)cQBW+8eWGR246Tb_+)JH@DS+W^g68W]H?57C?=0X)\_adRD;RO=a#Fg>bc5E
>-\eK+4(Q63\N.bG638[[DDP\A\5^W<ZD7QeK,()-O1_D>>7FBMCG#&=C?g)R6K&
WMcc3>#IZCVfY[c^ef:QX=L#[P?TWSWB56^;E/TR>0=+g&E^4D<(O[Dc8R3C2ZWZ
HQATef30>fWSJX3O<.g7b8IDG#8GM.KB+ZZU,ZW3Q<dY0<89SV1XK]#:/c7,ee]O
+]=J>UWJ3M&f^ZV7BKZ@Kc3[0)MMODI7Z@RBf,PO.;DWGbT@Y>)4g(@e8M@R^d/3
TCIbQ0?9HT:.>8M?Ub79];5<32UE4.ZWC4f4_1LD)U[RgL5T3)(PM3eYfDX4MPbD
K]>AVWLDAX9&>^g?XdDbPcR8]LQP,Hd9a[W?<-?FOWXIP+Bg[?1MFYd>:]3X&(P,
G(D?A&+:0V)(<c4NE65\7Dd7I]a<W_0XFId6TLV:RDNgP:]=XGQ]agHC_G)754bb
DASVTMPT[<_>D9XDFQ#]ZD]S/g&Qg>C+NX6V.P4?5fO6<GY]K;Zc06\c^^N:@6=&
+?QRJYQ,_8AT]96J9YE8QJd>^8@<BE+)\R]FJ#AZ?c.a>aaeE]=4OHbZ3O8VcYc/
GVK^dQH@cS#/N1MgdS54AJCc-S/VW\7@E#+XdHf(ZUVg>FF+T5&+U:(?:G6QTg?3
ba(Z]6T[0VH@XYKdF7>&H582,GHg1P86cYON@TG&D70FEQIE:MN(ffL>9S_]<&_5
;:#g^S55,+F);08+-A4FR0ERRcQVCe;;245]6#J)Q:=8,_MA_3RHC1<JNK#7cGYO
;9-ROZ_Vc.9<&QVI+ge,Y04],?PTQFC:L+1,489)D8,>>(NY;R^QHC55/g+,8<HU
FggXOLF,,&E]Z&U]LA-3W\5B\?Y5RS3Sa@]0C?V=IE5fO.->Cd,g)MDIG_cY[FUX
1ed1<PXL1=5U<<g_F[:FYQWcD1M39R]dI6L5R=);BKcVQ:2a^fWP^QN.3?BaHV;X
F,KIGG1MRU&5d24I(M,LaT&-YA>?)O<S?\g]:F_=>L#_;B@O8N08g1?;G_>c,:]b
8)Q001OL5A0,POG.@Z^I[W^E0:OfW2K#=?8GK(0@YXL]Y(W3\<]PR=UV)L;^3DdV
N<PIg>,+UQOeTBM4XA1Tf-RR9cF\\,<FMUXTgWF:8]J7D48bQJFRY#U]9A,SZWZY
Ra0E0HL+b/5fB2&E:K410@U70@OcGcA#EgPUOJ;&=V/O&b>0#(^a918J@65e9)XF
2?8#;DJ&UHB02e-+-R8;edYc1DOIK6D,9OVQ@F-b7>^ISE@11I2Q0XS__8[^eP<&
.1WA/GR&:J5dF0KNSca0af0aa?)<X-4;?T^<-dHIPQ3^@^@N0EA<M/&F-E@a?@_-
XT1?UW[g,LW9A0<>->JVW8JDPQcB8?&8?IXcY-Q(Y_Q12_SQGC6,QEZ7Qf+2[=;5
8@<+Jc0bIJY1-;FP=4@#.a5[7D>Ub/7fdaF116ff0/=]&eP:X.cCR6b<A):?&([Y
AIeF>&?&3OTV3+9?L6MLB]bV/5ggeU2]:(GM?3IH)g_<:F0=?SSGFeR3QW6?U9-?
Vf\(9S8SV[XD+^E&Cg]WGX2Z&,X&;(9[1^+9BS6XBNbd>5&&P\#8D:_NN9Q@[g-c
EW6MF.b4eg6C201gJeY+Mc>-/D[f&T.WP8?,\e4M-^?\BX@TENE;3fY3.W5..@S\
->R>Xb.6KAX.C-M#_5fb=#?FU:D#@Md93c]_Y1B13=F\VF<&bedYY+fY32BO^2BF
=Y0?aS\@I[d99)-/EO->)eMdfa>=5E,?^W??KU^T]_I3cb9Wd-af7gEeL]M4HQSN
=VYO]&C5a3-1K1OafT;)6:3^T[WQgJffBTT??X9S[1]+a(gAMe^Id;_O9#TT&R5S
ZJS8<D23E\V#,(<N6=Nea9)6&?REaC347POVVYKUX+;eV-7^9/2gSDD22]\N]F(M
<>YNTE_2=@Ig##ONPCIM3dU&=6<ZNg>;>T5)1:&e0^K&5PWX-=C,S&MV76NN\>M0
O4VQfZK_(Ef]VeEMZE9L<T&K@6VL4=00+cO2N98>D<a[:B-/,e+c;EY^R2+f_#93
2_gLTMSEJ)d0N=[)c2]e5YB3RHaVXO\_eRBGU#Q1D:IVQePZ_=WK[5Ee6+Qc:32G
RU57X[86M;,aSU7g#VDeRXFN]J=BE7:Ja;NH=,]d047c;gUW#4D@J#S6<b3D&e)C
?e(=F9a]4/Dd\P.FD)HF]D#7O,6]^<NbS(eg98Z.YB5;gLTTRC\PXb<3EKXZE2Jf
0.?P0C7W0J<P3@]Z5V&.#ZGIe&.YG63:DS)R_M:[KNf4Xf^:]EI6A8#gbV5H1aL)
WYeDHe+=TNEL@T&^fa-\63d2aVJP)D>R0P_<VfDUB].J7.-;V(]H@4-]a/a0:MO]
^DM;P+=4W+WDH-=I(8c[7-K&fU,g;&>S/SfL8U9LHIE-[Q8Z5a;g\1:d4?1_?Hb^
XK()LBB,Re_WS&V0g(b0c[37<7,Fd0UD_X.e6(I9VL9_Q^9K&e6,S8R]Z=</^EX8
\=DR2DJ,#(G5ZXMcC[.M.90C]HV7?bJ9K<MTO_9^XY<EBGG_]F=?G\fS\dQ-/GZU
R_&)-->8a6?#+[2ZC[_3#:_24XH^D(Q/CKZ9B)B==[<7_afbgd_MW33<TVXT9#2_
2HC:Y6C;I<X=Hc36b4H]-TZF2?@Of^+3^+ZC,T].LMU]+9&PeJWe]^09[4UH7[UG
eZ,]0_CY&;5T4[38+a2Eb2?DF0Q,-^MWQ>B/&7T&KQLdIGPA?e.ZUEVF5;Z#Y\0\
D]#?BIL_Y2;4eKb7@CI^7CO]85N686I_afSCLJPe]365#@<4UAO\\&4-)WfTD;XQ
E55?HV<)VIFL#T4YG_?(]d-G5/[+HBEL@(cA7&D,K[)2#CcSJP=8_^:Tfg/[U400
9=3?_,P^@g4YU/&BUSZYC?5b_fI#\]aHT:OKCdVC^IVU<WAWP?1Q1Q;H<OE)1@gN
QQU>\4P2Pc_a+>SPI:<YG+c5(UW],dU40K<T\N;2)/T2B-04>(RTYM4KVXF/B[\)
<61;&ODW&6,;?;>K1a3,#M#<6I;EaO=U55;_^@#B\KAGW@F<>]R&T9;5_O;fO:G&
EUKJ@3b+)1BKCJ8NCFCV5<&Q;-/aS[BdE>DL;TYe+&<8d0cO4NRF>gOAW.BZa+^B
UN.(1Z19cb.U\aN2(IH.IM?MF-NDCKA/>W<BK\b^.,0.F\Kg-d=R1RM>FdL[;cH(
g@+BE26+.T9&YT[O9X\3G0(3.KPPG)a?SEPNJ72LfEEOAWN>R1&7.(;L&efLEY)\
4\H\AVBbSMT\Ve@Y2@QP>@EFJ-(bXV@G4XQ0L-)M[gFI_\S:2?N^_+?a#D4GF?^Q
.@PbK&2+=B<?Wb\=DX,VGfaSY.4UFF]^5JA^\[HI27F<b2E5V?8V5/NY84?ROB,5
&V7=QFS=)J_4VdVI:EWNM-fT@cD#0C.F1#GO=g8.::&)Pfb2@Q+IFdT30f_B^1<Y
2?a)fBKDH,H895C44[3I]@,a,V4=aB;M.)g#Ze7#[5L.E.Zf?D2&E.O)@-]L7dfS
4+D^T^.A4A7OV]gCeB.2JIBTYL0GfMR)PZ_Sd>f.e?D^1g?IAB?+WURF-Q+.<\A)
DD;VW=>)f3>;-Q85b0?6\:D@#1eW63>bQa2gd#\0+6b-K3Vg:#Z_,Q+-1&KKJf]O
MO8]F,bU?aX<1,;^V/33Rd#e4X9VYb4ZH_@PR7=X6TbNZX>+gRTKQCc0./g2:PA#
C/NI)^F<,]#U-Kd^3CbIPMdR9WX-+XdFXR(3Y6K+0HfC<G:38IO_fLU=YFL1+=B3
PG#O>/96<=+)g0<.LDM,_2_eO8W[0Nd;XC>aFWddN#:>P[@=[^#MX\0]0(a4FXK6
G/5K+0\7e=(9U3MWe/5SeF4X08L(DQ^?-EB?c&H64LH)&++QZ>W8<T&/2XQ]e_]Y
Q-/5a-9e.>7g//g-2U@LM.KR(8J=a=^YRd&_^R7<gCbCN&HPI.W0gA1D@H[c\FdZ
).NC3HTNOL2S6P0I9fF,d<3fP0gX(A(-][Qb98XW3M:I5^cR:4c0O/@.0(TCV>5K
BZI9;-aK^SfNDQO2[B5/Q-R8+F-./V=FI;aYSCdgWf>ee:ZWP_(aSQ@:@]F&SgC-
E1]K,N-.EEL?D>8cQ]8Jf+EI.2AVBfAK\)-GB9@WYaJ_d.2<G(a9(_#5<PT2:?ZQ
)-,IbW3E^RQ<+-S;bTQY[f0@((ZO\C8109D?TE]U9]cg;O@V18Lf@HSfR:gMSg3J
V):@N+3;Ma-I4@<?M?Z?9[Q8MNZ1H&ZW5RA>7R>RFCZE>MM,HPX\UU/]ME-3fFLc
Z_4[NUE]6g)D;OQ;^f)gPKA5@\ZZRKe,J_6PWdWe-KCd;II4.I6\[I^FYgc<\-L0
1(Qe?MGH;UAV0:Wa@1+7H:9?4S0BDC8U#aO=/fXF^C/IAV>Tcc]&d#N[c<c^f&2@
7X/G_MI>&K+a/,GCW12G;R<gANP9BD0].LaOM<O#;VB+a0dK@-/(WS1Z-O,JFJI#
;e[J]Q/,NLR?L^+^G/?4BGH7E,NHOLbGg8PEcgXT0NXV>\VYJHZ3OWOLL?M8DH?0
1NF)W/CRHNgdI9VPI0/PUTeA2Y>,:+NYb;5U(#7#IUP40^8\8J[,\.UW7SYSD]]Y
P^ecPGYgP=UU-.4]L7RaU6-LUY7ZS86fM;dKXY3+AP3J>_S=)W@)_d/]&g\Ned[E
@#aUQE>QZALa#8@YPFN670RQ9L?E>B6;;BfZF=P@aT-VVGT=d-]bI#76Ed[:9B=f
D;?0a:gS?X8UCbTC]T_5JEJ^6N#Q,Yg4.REc_FA[S&<(C6cQB2_^.fF5J6UI@d33
J<\G)a(SBE)]1e4cV>O_,::\FAaK8I@P?UXg5)2?R<Z@0-#XW8+B6]_7DeR@72E.
\T=AgD\X9,XJ933EYDQJ<_Z+\1?_MBc1N[b-g@&=RRg,:b#85_F_@&0^U00A-^2W
DR0;CNQ4B-P3/Y[J7?gVdSEMAQXPe9e+N4<LI8#@)_b@,O]ae2HP]Ob\N/1:C3),
JC9B,baMLb#CBEAC6=(+,cde@H16=G:-LKS6B3PbPd2[+I>B[76fY<3(Z00[c1A=
YX[ObA9L[481dX=\S[^0]4Qg6^_S1-OENR7E,@Fc^EFA0I-,gWNHfW7K><^#&;<3
@c(]5^=DLTFZPVNc[OW)<S^(@6T/2<9>VD;S5>aMLC5[XQ_\8W,g<SfPM\4:P:8#
?K63C/&X;3W)(a7M)@>O),f@H^HE?H_M514CSOb&KC,b)TCGM^CN=>A<M9SN?#]R
HJ4U@^[QN6PKS#K0PeZTHL/W<(5U72EY._,AIIYV63.7J+.XDC]]S9/[K).V0fQL
.+eQT_&A&FT(#&N<H6?cK3XgU3CQ<-IcA>-H/ELeV=P3,FL44=[X&],W250B<9?g
+)57G5M4NSRO.1<>J@21@HCJTP=bJDQ+Vb,V)H#<F[BT-XZPd9@I8DfZ,+g.I;NE
Qf>K[KSR]f9^Q6(B=V4A#^0M1@#fT6>^,_ZaD59S@G/KE)e-Ge8Z9+e+_D4G9f?9
V:bVCcG[I97Za>Y&b[ZZf>]M^<]3L33/Q^X=@+,eA\d][X@=@gC>/H8?fL<?K9dG
S74g6P;eVK^F#U^-BZ^XZHA9Z&=6eM^]S\\YOeL/V9S[@_EZEX.P]bD\>6LFU?[R
NUT2;BYF?J[8c)U-).7YS8L.GY/T#M)V9]M@6EQg&D3DcW39X+G\<R7\3dF@\<NP
27&LS^cK]H=EU9?\gTG-?FOa)GU(#@W-AVLd_PCa\&R3fIY:NQR19YLgC-gSHebR
;a(#R73W\[\A+QGI1L7<4Bd]\bMC3)@4ZJbC5[_##Q\,JYS;-.K:&C+4dMb>\B04
.],c0M[];7PgNe2&S@GB9KNWSO=25;<@9V<gBRf&2/P=aM#/aH(ALP6<LW543OK@
4MccP24IX-Mg\]BQGaK^PH(fUPHU;4dBe5MR#GB7S0d[FOfbFO:,^3@ZN2&=>a/0
-1a6SDC0UC7-Q]2:/D37X:D;O-b[WX)74J2Oc/1O.U>#0NE;RJJQ4\aQ4HG8+>dA
.9+bbFAUSIGe@0Z:6OaK@E\]eVEe:8fF<5,>[)ZC#eN(F.9?L=]+^T,SB5KFVK6@
dSW-P1N>gNIPbea4TE(d4V.6d.IMdEYY->M_Gg3<&)_GeKCeGL.F&NHWKT=DD=_;
F+EB0CG[0V5+MMKTJ3dfH3AF(9BSTHH\>H]OUgFR=GC9O2K?dfRZNCNU]M)JWMbP
0I63,d2)1(c;83382D_M)cDXP3^aFM:ENMA/Z[9X[NXCQ&D-S=8:3@E#d2]A22S9
<,GBFT>Tb.dS^;_W\I+c;5gL2c])3IdDYNU?^3QTDGa2XV]YX,I=XFNa#4_L+I4R
dVT6)6AdT^S(ZKUJWG;V8^B0_>@ATY;g?8BF\AeM(+&MSOSWd&Q;5;WD(V<2+]2W
2.29>>S,IOWS__G?OP65NW?FZGG_NdXN9HOTbWE^<;EA8B(?G7,INR5+N]+C^O(Q
(b7A34;MO,Od,L0\CZ<3U-\O#Y:]2UI?J@)=>4N.&5CGGd-;FbOCa;K&N^2S]9&f
NV71AI4/fCYRVZ(/7/;dG/aH>VT=:OJEb(cQ0ZUFI>6;bC@1/FR:;UaXL16c5YB^
IcaL8[QNg&UBgZ#Y40I[\JRO_:D\=BO6KaUagF1I&3(eTDdR/>c?7Fe<RXW+d1U]
EBI)2<>=\#SCaK>\f088)U\SNKcb-=#].bECe)g7:N&V,H)07AZS/GDQbNHTL>M^
N=6=.&e(98+PZN7\ND8R4<.23\fTZI<gQ4E75)SS,IY_,LHJ6H8.F:aa3bMHb65c
>[E_f)+f&^3b8YbLX\70>S_1G_FI9NA),YLSXf9TaWE>VJ<(d=QBEgZ]4e\1ZL3)
O?\18:5E.;]/KALB1F@0NBLTJ2bC:?G4R61[:Q+<_.A78-Ug(XLU898SJPZP=]-0
IPVW4b&1#2c+OF1HEOMGc_BN.R;fDEQ<6^LcQ(USU)Sc1<L-2:ME[(bX7Z3aNDN+
?Za79\UYW/3De7PIcAH4ROd3Y5N^-(f3V62_>?fZ4,JbWaX?:b[W_CGH-)&4V-87
,M,K=8?SVS&TQ=A:]18\dH)<2CTTI<?I[:R.=FJ;IQUQ3TO8U[1Q<bbY]R_^[>FX
B<-(<3D]DRb0=GXN(X6UXNId\#<+(]YdBV-.=I.#)f9TEA_HILJ[54c40)H,E7+7
#<T9d>g5B7ebOYK+AMG(5TDRb8\H860VTBI0L.cI-ddBS#aG#W^#5Ce.^3Qdd.fN
Q.<.[V(5K:HT)VPX_@\TT0LG=a-<d)-Kf7,).17CJ[SQ^e8MY]8BBI,]+_a,D7+e
3<VeU?@6@\d\[5e1fQQ@B&U-Y+6(^UKN.c+3Ac;4)7SAcfe@f;->)_eWS/Y+T7e?
(V3)NVVR)[0aae4TKUBO;@4B8=:GN1,/VK+8=?b_&B<1R/S9[#E(d&b^B@FW^Wd4
fS?,b1U?=5.#8O5F[SRF,H,?bV<YYY+SJ5&fDB:.<[TAT<#7NSd-289;/acU-I\O
\E.^^&5]._@H=+B_37J@YODYcW(f7K@M-9R\/>-dbgVfMW7R3I2cM78&\Cg^-UbO
0BMD\^0HHU#bdF^c#J]A.Z+/c^N>fc1>M>0eL\&Q2fA:9b\1O/-Kc40HN^GQM,&L
f4?P+,HfeWR:\RANaN;CE-b4(_P,SDXd@D=g_..b_ef2@[Fg^+SB>;DN9^FL8X,H
XL]@>N[Z\^J3@0]+<V^ELL<?fNI&PY5\0d?7C+]R-CR?UE+@b;OSeZ_-G-Yg.KaX
#OAN#5UCNS&W\:.1)[1Jbe276O&25W=a(V,XWTG0,WGDIJ#:f/[eZ?>#1QVe,4L&
?RA_<aXe6J+efMS3&+dL+;QY,V[+)E-PT))?eS.-dVOGD\OZdG?]WHY-O>1\//HI
(/>_C5#<=SgZ;=.fB&2_CPgf540?7987agR\>C\3=,NA+,RRY;YOZL4#[PgH6C,9
@58,2RPMgAA7E#5eJDH7d/7#GW972/7DFe#NCXZ=IY44Ug@?;[^2M[DF8>-6#AbU
EW-<[b/E1D1UJ:,\003fcU1SX+F\4bf45,THdS#cPf#QEH<^P>SY,#^)P<Xa=JW]
T2/?-7Y@KLHTJR+84dBR,eVZUI<Q]7ISeP2Zdg7c(3[KE.+U[5LI/3@LL=FMdEd;
&4^(Agc9/U>:_O\PKeHbG=Q=,\Kc)bA#WR(d=.L7DO-EE260:g8ec/XV=>7IIDcD
4.V<HUIR@>9TJN./X[.P@N83#>K,Mg,VQL&>_a1R]B9DI0Y-UbM_9Ja;caA&N#d\
/We:LSH[3:77dYC5R1632&Z3BcMN=)+L,5U=Ig5\9S99T^);dFgQ-eJB6^L9,T6Q
WBW+_ARX[Q2<)C8W]@&VgLTQ_HJ2EB82M2S.>&PV:;612e2<W>MTDQ^KUNb:I322
(7H5QYP99fD#PZ>X_GIcO&I9#;<G<_UW[I.IG#^]C>O0bVf5VHU^>(@=+8a^_XRD
DC42H2c5XSI8]&1^\@Wb?56P;MeO(S6BI-XCQV9;26:21fLS;S-I24f<U0S3)JLW
<&ZJ8)+02+:D:FPg4-<8ede)eXR0N<<)I6U<4@?H>2E#H?VY=4Fg#_X-Hb@;9(&+
R[5KfEAgDLWX:A4DE3=7R&KR+HcUBA#fI]BO=X]+>+,GYCXaN[P-;W>@=&??87L=
M-TU-):MLDKHLUVf,F67F:B=4MZXTH(&]^9AL]3/WG,]dF06d.)ERIRATS4P^A96
OQ1MEgW<UNddH/)+g+gW@93WEQ9L/60<#3S-f/a30.g1-eWXP^EI_HN=Q+QF]_2N
=\QUJ4R+(gC)UP.U=Zg(--gA5RAEJJ66BDO_[\d5BW]cF/8E)3SZfO:B5IQ9?bR:
8JVE7O[JWZ#6,&ZF]gX+eT05O):KM1RD<0@+EJf/DC+E2K79gWOF6K=NHO;]OLH;
/g2_G-<Gb@;3[^6R[;;15O:9(@H\L#[T@[#e,JR_UVJAHgU;18_S(^H8+/,Lb2<Z
SAF4@1U\abRQHGU+>]S>3UeFM@3:fff_[ZA(g8\WCSXQ3b0/]:+[g2>#64L2=HUA
@@L+#dH:=MN40CC.Z(MIX/@+(KRI8]4DU51S6FafbA:bDAKYEON7ZHK^]L^Fa8#g
V&@D.P0R;7:VTXE0HHUW=JF\gR,Y=.Md84JM3BJ:G69U:B@ZMEF?F72d0ga#(,VC
e&P3/JDWW7:#0:c02;IB3S-V6/BYCP4PA#.L::]N;0BVb&PK.ebAF;#GaEW^gNT?
.XfR2+)A#,_>DQI)O6Q,(-=5\HR2=ANe)0I8K7@R8YEK0(2:fE948<TMBOLO,B\b
a>G[,/WNb7=G6A>AS0E&<S]HQe:96J--?47Z<+;D5c;94^aUc/WbLf2[IS2R09C(
Ia5;)KRgCJdCX;?GJJ_KPB9^)bA7,]6Y+b7OEVC]_cMM8;L:NO8/Z29c[DMDd-aJ
K509,EA0V;EQ/FT>W^IW3]2[\I>6@7:N@@NS_AB?@;CK(.0a3e:ee]E>Q]eY2SPO
MBaUX9DeU5HGJPLG\^?C;2(#D6C6gDPI;^gQZ@#Tg-WgP@DAgWW>=Q^KBT_DUUS^
9QK68(,B9gE]fccG:J_&?<bU3=7g0/<..bJ??X\ac&IT#^d>9H9)I3)_<AKc=YSU
>V,3J+WN@TSL.@?5^996-R+UI0)T[_L>/T,2c98#VNg<_=JK7DOZa/I_P99/c?Vc
b.S7CPF.Z2N72=WI\DaY6-.W]6LUY5^.H1>V\gcg>EU<\?=@9a1^97E&Ic;51WF-
cLMD/B0NO[[4<#[&ZRX)R98BJ(\CL0RA0H,QdeS-J8c.<cLS9a/BB);T^eA+L]>K
36Pb6QUC8G.-.F2)d/9FOf8DO3LgJ1:3V_T/T>UcfUY+eJL.eRTb0OEV(.Md[a,d
61QN(:.dWe=).E.K]IeZ:I->2AcR@dfI5fVPC>a42>(1a@_K763&]K:9XP7)g/QS
-V_5P]3-H<G_ABJ:_?a<dVd.3ZI;aQO,?D@EX42SX9=HYTLC1-,[(e?04GO#af/R
;c@-eeAQ^1;?bQ(26@EN<3Z:GNH&U[?2XDOeKE8IaIY/^9QZfbUUeO\]V=@O?VJ7
;5(VG/^9]CBX-_3+X/,G)FTQ^bgC&Jd>(c:)V)cZNG]5IQV.VM.2b@0)8?YXQ9c\
48CKQdUGdR?@HF9[;_EL3728)TfKFNQ;?<f65g#d,GOZMf7e2f\gMd(AeNUAT0V8
CMX-,1d/,KgPP,+-2N7H#?+Gf6N+bX7>d3181X2XS?P]YU8RE&_/K;9+8QJ-8(Kb
]XI#_&_KZH[(7V?Bd3;2cJL<5I(&7VQUJcX@TU<-ZaQF;0=21N^bI=Q1G.NV\@K3
aB?NTE]>BfX51JL<VT<J1X5O17:-H?8f-?JYCf/7bLZ1=)AS@FAP[J+.-Va-IL9:
HG#3(gHT>)MIANX-+]g5J4:[JM9BC&#0D=)/5/TD)?<2ZU9W6Z;]TH[G==N1I@<-
_[&+7SQOdJ6AbJWZ4dEfcC#2+FM,JBe9K&dU,EFC.BD=RCFP.a-9<7MBE(Qb:V]]
c8MZJ)-Wdg&\WKP(Gg-?D#PE38M(P_BLV>c8MBgZc3:.=0Wc7;.(Ad4-a-(0(K;T
DI70BO4[-bBZ_Y0TgZ1N.)HbCT;=WP5&&>gDR[W<gVeccE(<MYA?0NULFI/Z@a8T
JDFMcdCNCYP\(,8#/TM2_4P,f1<DLC_F2E?g0-IY-S=EX@0U:8+PeK0CCW/3=VL/
MEX3Fg:ZF[)Q1aJg([+Od6?-f8bY=\_1D,>V4&HM=Ve+BX/Y:43Lg).LDKX(+dR\
9D^AQ(+E0Yg3D4\0D:>dJ#H.;\ELU-ZYYV@OG:cU8cdFE(afb0G7:#D^;E@G<?VD
E>+KW61/HMKC2IS,9\;.;W<NDW+3PB6:0/d_U=:]Ud1e:.[3(FRC)J6dPENdg@10
-Q;[O4J8ZMF5[DLNY>44gM5:Y9GTC5#RNVA=CK;D?[0(#58+aBET2<;B)--[<+88
21B#7F7(PZ)(b.VKB;&f^@?:+NT;W0gF(bYF<;B4Va/4Hc__<H7g:F8Xe@:a;BZ/
?GV5D5NeREN&7-CU&[LG:#Nf.1F[9bdg]EV_<:+d3?c>1X)3<34-Y^>-UH(XY.8;
#L3_Md)a7E9Q[1\8ETeE0YfTg8@Pe>B\(9PG[8C5[PN((-CX(]/)@[d(NEDJG8EW
HGC\X=;[e=(QVY8:?I>gR5KP.F7B4SRWD-g_(MH407PK2cO5YAOVNSN;,gd#Pd;0
15:]WRUI2VA_H2-a.Df;@_7@CJ9,OOG>]eVd)CA1a)Y<5+5;M=)UC4F1J.g1^CB1
a4[N4/Jf7VN6:dePT@cTK-f@^^_;CAMb?Z)D1T]B(G^=,8;;]8)1De92@LHdR=;6
CD#0B#c-Q+C9V&=;J.c&g#]6Ug)BXLQ<2Fb:G,_WN3&&B,a:KD]3f1^R)6UeEMXG
0NY]TT>J,+O6:8T[:79cENPR&BCd/+F#EAAYDF_=^TUPfNPJX:[5K9BJP]Y\aIH8
QdA_]#1CT2OSWU-gT-)?P\C^A@RF\M/F3@-I;42C:cDdNT@^0I#6]2S_\LK=220R
9;8JGGGF>KX3U5,-M#B^B:<T,LZ9LY_4X4;O?cIA66.XQK5TGK5TX#&g&gVF]H\@
6bCFN11^;5]T#9Ag98]9@SMC<[5S>K0&0Dg.4ZP_NC^_7GXQcH5AW<QcR\8eT]F-
EYc+GAMcQYO9X;_L:F(S#f<Xg23/-/U\g?&H)<X&&]&>Oa73FYLaR?J3g/>0L15T
T5<=g:-BN0>ggf517W(]RW,D@;RTc:92<[THfGbF?4b@=H03:F2g+fTSXdWd[cFK
89YL.F6)HK,3UJ-8/9&MM9F:?G1)9T<?GI_X^_]K/D.7M5Pb4FCY-2-MSH\?R83,
B;c0.=PE].aQN/JXcZ@DN3?A##,_Q-QH3c=<2/b539&R^C^\QZE6&aW;VK<<4/a.
ERX22V/6\28ZcAO-J\9(]DLGWH_]b6:CYD[ZHP[XbL05EGVe[T4&UJZgYB&TM:g@
QGKEXQ./+TTXe)-[12[aY9RU1BNG5]3=GY.,TQ>a]M6FQOEM0S.U<\YIQ-ZJNS1D
f<P)a3\0(aSS[\47?:CBO/=_.WD^Sf-?L;2P@OO:^-JQP^f^/a-G-(IEO0UbG,?d
0+>U>.aCRG3g;(SYW(X&PdO,S)A,,3&_cQ>T0MYS)Bg,YZW\ARK+]+c5bCZC\QY4
2HD,8(+8.TKKZ1&SFDL=c;_I_8UA+#LZ4e0:4P;]I-67@-CP9Q>X\H-NNET,38:E
f</1D^(L.#P+WDADc)R.QRH0H)-Q&:\+;gY+38_e)F]ER<[+1&g6g8c[J5ZdVH@6
4?Xc^fYb:2DK=W3Z;@G.WdB7K8KW+SU,dA?6F]14a?9M+X+TPRD14+Ge0YfOW/Ic
fFfDG2=^<?H,G;Qg.9c<VQ3IB#[9#dK8DFW1(K;6C,=;-b1)KFHP;XV^8_Q/+O@a
Xb,HEf90+]FVCeAdSTb=c&gS;D+;2S)3(\EG4b0Dc6T->;Y0N:&4GY@SF:O;C.O3
bAFVT(G1([?KS@;7:;10LCSdXN-T/&9CE+S=ZS13#ZEM,:F?RO3X_c6RO.J\fB5g
66Tga(A7-ggJP]bHaR@FVPM<#EAUPF(WQQU+YPI?.F\7;BC&<Ggf+]G(cB2^Bb9#
S]5V]J:47f,[T/a/R\&ff(b,P6d=5JM=)\b=A<OSBRUa4dY+HLIc2aQX&Y528W+(
?>\+<W)c&L_<GF0..+HZ;S31.FFJ9g5-8a>/@M_9BQ4)9;I1CK&:.AY9C9W8[g_b
G>A8VQG5[(bG?(YPE7JLE\;d^YZ_QLRE&[W=Q(AB)Z:QK)b)0SLY[XKb[U0C4J_<
G:[#Z)^A0-2LQA:6Y@8-]M[Q,91^OM/4\cVTW.GI8BZZ[[@ZIaW37\5:?8G\RMYd
U5I8PB#-/(/V(\DcVUM^eXOUT+GCR1^I0GNV/]a-D#4@[WXILe4/f6DU#:[:cNUA
Sc-9c;egPBCc2YZ;4f6QL>,K?2^7<+]QIa&cS]->&6N/D?4+_Tdg8P:D6L#X2)D^
R:MeJ6f^RZ.#4AAIAQDgH=C5+1H75(9J5L=Ue+.CfS+<)5KMP(O(DP48+9=XG04=
326A3[Y#HaJ(-_7;dP)62?[7&#bAE/H7f_NKTSRC7G4Qc(G5Z@H&2f26Kf;@QKdS
4NYXcV2gV9C?7LCV@EX>dV7YOD260bPZ(R<;TYI&ZF-d8=dBOfQ1I\f9?M<)>1/_
Xage[:H291,d61QYUD-YB\+4(1@50d/X?eIL+#(LRV#=>>3,9FI>K1A[,J=a.2B&
(YEBQb.\&OR8@D)6ECSa-TU6FCP8RB8+9PLH44U]1Q99bNK6JObgaTJ\#?)2XIZP
:T@bZGaXEJ.))7f2aKKWK6QdI3[CP/A0MVMS]T<[/5L>M;ga\WCLc[d5,/UFZdPA
WKSaUNB[L>7f(Za.>ZK@CS+31;T.])>&L7.Q;9d0KIUA5H65GMPb6g1#@FXLUY.=
H&N4Rc_:&&L:2<--LY+g<F@RBcTA:JbB^=P;g(@^]YJRD[4L5SV>PPRVCTQK3O?S
L#N<P9gEHR<T/,6>+XNPc((B0SK8F#;)U4T&dCB=\\2)GLAQ<c<D#^\=d42]RKcC
:OIGGeZVXI:7B:_GdK>@NXH9JV1]&KY0eM]-+\N7;T/GG(#GD\YQLJ,\2aZG<e+O
X#3H(dXTEYC,^JQS(WV>91F9VPg4<_7=U>bTe6bcXK=]ROV5-eNUOD_2<:ZYMSNK
1C[B]U(^DJ?=&JRY9YOD)RI#EB1cZUULJ3G+c0#G/GNe,S0]Ma5#@HR=QPQ&0+(F
Ge/ZVbOJJZfc7+W1VFWU;<R/R0YCQacU?UH]ab,#D\O3cPZZ3#3]08b10B^L-S4[
M)M_@6UMeVCaGQR2\>;3Q8+J-:L_14E..5(>M4bP^MG04Y6B<B&(2L.fMOBT.bCH
XW-Z&P@2JT>YCXH2c=I&NKF<&WAP##JR#g35R>5gVW.6P(<&F?T\^9<b66^U2Hf+
8:a@>4aW6O.Y.PS^9_aI<3]Za-,Q0LJS:/@U-RD=]bPV4.VA447f3L_.8I.\acfd
KU(>S>6?9\K[DIgY70W7M)7Gg[<^[6C1NI:=T0&gd.G5_a=[(.:a=BYN5K-LCBJ2
Aeg&FX1W5ea;KfQPQ>I>=4DELe2b&6JK\3KPRaU/EKW(5LORH.T0+\3>GAZCCZ_)
3_\CgZR:cPQN&P0d)WV,cMa46\:]7(Zd&<)O49dF2[fL14Ma;cgc-LOR<a&[aE/9
@7D<@2]<+YBJA7ee=XBJ7QV?Z]1SHV+YBdL/]\967<WG<K^X?WfN:68/Q76N(X,g
7ZQ7g(=b3_WbQ)6_5L2?7IP;0V&\W>+_ILOF=H\N9>Rg8e]L[_eS6)?45WBTT-b9
U1TBC++H^ZcIBXWd2)<7O=J5de?BYeU3;>)0Ge^U\b)aR(DaMYC;HNI,OEH)R_0Z
GA9G<AWg0U-5>AWa0)KOgUYPWTB)<O[ZCKQJ0C4TZR8ALO3caIa9)NH)HcB^gM0L
I_[7UHd@a)BV7\CT;&]SZGMECd.eGMdUc+c[,aO;-)gSR8DSeCJAOVfO,7ZJU)<8
UU486#fYB?0H>?/87]GK0^D?@Eg#B.B;-^)?\D<6bC#We#5EHEH4bE3CW^EUg[YX
ga84&^206YgM-S,,T63.Q;MX.:@Bd34_=G=KM0NU.QeHO(VV7NO9SM;Xc1f2,^6M
ZFd\;4RIWM?TE-\1.)BS1dH4H2B@=&R(YJ]4TP58@(D[UPOM7TA\_77ac/.#PPE1
dEBWH#g(;L>R2D#^#P]4JCD)=Ff_Qc[EM@e>7OC]G/X\9B;F^;,F>KNQE/ZKX,7O
eEIJ<7<gGY^NP^)9e,5HCQ\bCHH+X[e]IX;9>)<8:P&1T;c^DU6JWHc.410,-e)]
.Ig^@b^GLTCF<3DC3=K21/DFWHdJL+4CGb,@,?6=&0a/?.d90gaI/cFEXMA-[=Wf
[84PLRJEga<T0\_EB0])F+[N)4IJE4,X&dVZWdd[SRf[\D97bJ,V)E&]3faH;Od(
0-B>Kf>&UD;9>G=<LFZ0&<=f49a;@eH+IV4<2c)9]Qd)P2XM(f(S2aGTa>f^LBPa
SD/;\aX/=M+3(2N/DLW5c08+3eV;OPUebf(a-D6b08DPc#P/XF:HZ-OfB&_X2T<[
2dKE6;5C#>/D]S[/B_/&><&+^]Eg(J=MT)(d4&4@K&><b>3P16B_)S1OV#PEcC_C
#WMXC;(A8c7T-Z[SCVgNFZS(d<INYDD;,_^[dOI+/S=6e_A])=OZRG2Z\-G<&7;K
)5_C]b\W=;<@P-3:@/1YK8]W(91JSXa8(781>+ICP+R1@W1e]gM1NE9DCEF1/;4;
+7X8AI,Ee=T+&)b.M\)HV5c+6;DSXMY-HdfJJGA<#cV-_G>G,D?>OGaZCE8)cZLM
88KO_Q0.QgT+dZBXLU7g5ET(ISF;(].2ZKMKO1L9&7XcL)gTHX+>2e;:_=JZG@[+
bE&CJ^Z[K:6PP/D1]^Wf>FY\2gee+1dVARc]1/X&OEKXQ-@b?K<^5&&WBRKBa94#
>[@1.3(>;H297YOWb(G,[,1)W6^.\BXCG-A1<(WC&5agg013XdQO7e^.K#.:agde
?g@2ZC5N1g[H8Y8_VSN/baL:\0:-;-,ab==7-_QWNXA8B/a)&#S_9@?0YU<;^4O^
I=6Y\I>>M76LI5-,SaWQLI>\@bWN.F1F)3.NE=D\G9J=@MeO+9Q#,5-5W/#YFS2F
]4JL8+7SCQJO]-O99N2/7GPe#&,eMFf>SRIBVCd\.;f=V7]AbD0aM8LeB>DX_HaE
d;0YFaQ?+Ad;/<S&aR]-T7.,#.cY8UP4@UJA9R^@fO/5LEgWI<+g]N^RNA2M3fb&
JD921,7]=82YUWV:2cD4&ZGcRX,bf8I#H_5:K/d@?e\A()Bd>H_Hc&E0I=2Ydf+5
dSf291YbRH.G9f4GR0=e?VB;D>_F8V83F9bV7L>XX7F4T3A53a<bT,4Q1d4H4D,G
MDd6c.aM(&Waf>fMGX]K@ad>4V^0V#Q4^5;^3;_@>OWHab@N;1IL4MFe_K_-4-eX
BSAdW63/?J_5;W@RFd#5F0XV(E;VK2;NV-U:L1AF.HJb6.1I2E3KeE??H4>8XGM^
[M50+5\,d>)9c-R9SGeD#AT;]XZKMg;,B@F[Jdg8K?CU)>P0S=?7]a1,eAVS.^?E
6R5R7.Hg2=@-VEB-FD8PIFdTAS>:.BPJ2+4J+?O#UR;:^/FcWdJNd,NGB5)JUP87
]=0CL^D#4(B)=b-VH0LXM>0P-/QJ2P:CWCE3B=>Ug49(E]OYdN,F?Q3F=+.5@QR7
aa1ZKOb+g]a:Yb>:#-BD<TDWP+P;7E=5Ke\=[eVOCT9CI)=/DD.2>aKcH>YX/@,K
DL(7#A>g]46Z)&^0bJ8FDCFM?H;g8\Ra92eH5Q^&W_.8JB3]TX3]WWV)4M^g/&^)
0ZGH^?<YD;-FL87f_<^2[^&2LdC=OB.WHZ2OFSQR2V+d5]d.4g8&PE3<^US^Hd[?
RTNLU^\E8LWA3:54U^M#?DFGW]X.VG8N-)C1cXY[e/DeJ#94H/L][f],&7<7[Hg^
RFOe)dZ\C/W285b(e-J2GV^F9fU:KQcY9f3:/P77H-3].M=_;TFWM?Z)TJc3D0@5
bdT3;_MCHM&KP6;XNgZB)_(I1/>=L,IK2Y&AAY40QF^PA+FFG7WDH<e2c9@)Q])L
X8EG#P6ZX<\e7&g)We\>?=/LcA\ZVCH\@T6&4_63.-JMK3O>L?aMb:Y-P#=M#<Nb
DUSB=99^?>E<LZDAg6Y82We6-SRQ<fdBBKVVH0K#3EEB6&f.-+X\_YH&?,2C0BY<
@IMBR>X[b(^a[217edIS.BbLDJ8cWK??93g4(;CCF7,^eGWRI&BP^(=/?X7QT@&M
\cZ+P5eL0g:f&fQNaf/XdXN]NW9]>4^SP^--e<-\DLS(&:H>K_M@WILXCG3&FI3a
U[@0gFG#]DAP7Be/_6&+N-\[e2/]Za?LVE.RTb_?e\BP<2BdQ0gQ(=SM,M@UbHRE
f4TDY8&PG3>S17&,S4@4Z^bK53)KgZJg3S=6?=+96+H;b^=3LRXg8Q0(^M&[TT=O
UN>K>@CeLXYXJb[UZU_6:=N7AYb7EFKV@([(-KfQ]J7N@c[CI&V4W>QJP-#FgMED
5:c0X;TYQ@bV)B#V_)bTGH6S.7U;BObUWd^c&Q7?.B#gKcK+R;fUZ;Pd>L@3PF4S
YHQ<,V@@J2:?b]^UXUgL8U>,0]>@>_E]GD0XaN+IWKRgc#WQ83GNFfR@E7[M9\3H
[):\T&U]c#gH]3Nbe.D,Y>/K-:Q<U-9?C7JH,Tc,=U#Eb\M)XIOXVUX?YBaT8P8O
:F>dSR(>=FHbe[5&cHd.KTcGQ(^H2MA1X)J/Q:P&F/<67VUe2+LKL6XIN1D]<7BB
d>e=FVe:WI&0X/+Z97=a/>/gZ][N8RYbc.gNUN[F?WX#<e)-A9+gK#=0P#dYI&Nd
&,J(V[\,XZgBJ#@3P@IObUE2LK2Z,Y(Q8F&N.ELNc-d&Cc4@+(0Hc5(R.:?AZ[C_
+/[Z,d2CB4@7;NZ9W@[\bKPE5HB@e6JP03+JTQ[)#CV,OS@[)\cN1=OeW/]F.N)^
A(3JCYMAAOA++M;(V==&7Ca4N\<]+V&Z&9;8QA2G+T,V1KKS;b/bG5F@KJcP6)FL
B/\#=Y#E11O0ALMBSU2>6Mg)CM2/#.@2:bAW[E^)JGJbIL5GdK(CYK^+_?TZ@<&M
-\HU76[N0H1NRLa[W35F\XbJfPf5(bZOQafTD1_27FU^O3.f,TB#6b>c&K0PG.Z7
[;#EY-0ZMce,45b;X:8a?bD8#f8;_\OB\ceZ6=5fSS34OF98M&.LIFeSL3XIM/79
(?=3c;62<=^^JKIfI10.^DSNc+UNY]7A8I#F#9fT\[KJJ-0?]E/DM31GP6D<3QDR
#\TB@CW:K;Y-7@O[8[-@7fg&6L1T=8,39/6R>.:YZ,EUOGdZO4^XD@C7.0L>fI?/
;Z;Z)13K9ZA(W94&,E<8c9[+[::T[2+R2#QT+0S0F,ab)BF^IHNQF(I\JT<O?AJE
RfJ3Ja)GSLFfd_<1UB^9EV.CPMFdG+]6-AS@eL\3W.((-#-dW<B4<P=DSe1WVb/N
)IcTQVZf#d,_EGXfKN.E:9,9>I>,]R+)WWbRXC6@ISVLCZ:+@NN;<=eK<OC8.ccS
2DNXFD>ON@IPBP@5O[70KX4M3a/J8PW1TI9<Re[Z:;V1@39OFRFVE:aGPN<H+c/-
c1=L)SFLNc<KNXQQMO:3:07eN#4G>e2FEO?aI8TLd9NVgTH.]#8T9:22P]7M?WQ\
G+,T:^L:A<<^;R/dTd_K4TPHXJ<a,fPYX<OgLdA^eN-T@@>MH_\+e,=];.Q+D;Gb
L3BF&@8UM-I@fe_B^_b+<@UdBIV4:R@_O)+XfCL4cP846/J-UTF^OL:aNff9GeO=
=XT.8#19L,6c?HI<ZU_A)ZF2cb6Ld>(ZI8\4V/SA>0DNX9FHXI#f9IJ-2&\WSLO6
@;dX-d/M6=+N#cUMcXg(@/(0>baa:Y\L0&ac#Sd#RNB;AgQ#A=9e2>gY9:cR/?M-
-Y:<]IP86&eY_=/O/1-^08,FQ+,AI@9Ee)=cE721HTBa)WV\g+4b81]FNHC9XD_a
9c@D\ec0ML>&@dIca8LPC>;VU(W\;3<RH=:DDZ1+\8OG@5_5DGO+]\J?^0.b15>.
)RZ&<S8K0.V<S)dZ-S?dP3)>MN9e\[eF-;D;@LF5^1):3>O5EO#^(D:G=&NJYZ:[
6G#:6OX/^4_BF=aIbAIgBU)>L77Bb#NE8^f3[a[^[4X(R?6@(A-D)RKIJ1_@@7<:
0<(\)CP1KXY2#ZUcJY(DN>,@4J9RA(7VI[Ib<WLC>gDH#CMMaLa@JKV-dZ0:XK,W
bZD56Fc-=@&7A&cSC=SFNW4SP&>/3+a@-I-f61gG,H+HcON9Ke0PX)81ET25<\Za
&&XRHeY:O8\,O?+ZZ;R76I>@1V9Peaf]Y(1P?cY+UgP-E)[VB9<e5C4I\PZ5EDa)
Wa@JN6a17Z-AFabR<V@cW3ZMG/S4XQ6WLF3fS.g57Q7ca/\g,7A3WI3T0eZ/4WgM
/JTA+bPOI&9C7XH.bYF).8WZP)Y/TG\J4+.g&736.GWUcZ=XFN-<?(HY<1I0^RG?
4fMBb@.G:W>WgCIf,559g_]Rf;LUGGGREM+3g?OR;CT]Ub-V/d4;/TL+CF6NR9LW
J/78-NCO4\P^c\5[MPgg)-f_[KMFMG7@GeCf2:W.KJdS=>>+L>=W-Nd_6]DIWUBU
IdD>?VJT^-a]0)DT792(XTLYR3GQ7Ed+SY+>NR]BMK-TR-]YSD+>U41>/EDP-UKC
DBgeRb7?2&(UXRf4SYc1/FB#\H3<PH@(gSGW/&K4WE&NB)1J[H:9cgW:T][(EOI@
/1S1,91]#H3YKWV0G=]\9XNL1SPS9#N=8]e_Jc_4bR-M5A<\R+?M.&P-+1(?JV+V
G;GR5,-KN\KfSU-4DbW8UDO4>MRNJCO5JXbQ5]8P3aMPTP15H?A0IH8ge:gG>#8#
^5V:8\)[d&/Y<Ja<J91,7==LcRe&:62V=5(4337d=V[gY1=ONY_##23;Y2G)M\;5
7W?Fb&^+-NbL]0H0Bb#5^5>e1bE+J.PF1dY>[Z+fOZM28EgYRb9>X>T1J;gBO0@(
0<D9f#K,].D)7=PaL.,J1aJMGYf?eDBY.>6TZ??AbT&DG,WD]:+E.J0FZZb5ZAKU
205H^Y0.[C1A>Gg@P6GP]2WVe-bC0dRV(g3eMB0K@71R]3AegLWf_KCfK,7NE6,d
N6U=R/-[Yd37CUHcILN[-)gX=6Yc^][NV(@\4aKJgH#08dTf[^ELP=e8UQI4;Z\g
(?IZEKP--C&N.-:O3_5J;eE5V0WKUAIX]S=c)cRQY[,\a#]BDGZ4,J-E6LC<2WNe
,G)Lc8#O0^3,E;8[V1\@>[C<E.[(YeI<JU1Y5T#cGJ68Y(/7e\#+@bAG=eZg,<bG
E5=,9W;dgU^VV7IN[.)#Y7P.3d_M#XF=S3=VT(:<UX_(@M1=<<@16X][Q-,-2&PH
^\QHPAZI)PeB[92A;34G0_3C1,.8V[LK.a0;eI/).?6ZZ\a)X3C27[PbO9JWVCKb
F#D6@0F_:[KX1Z,?1\\OGBW5+?.]<,?c98R.bE;/4=CXb.ODFgLNLbY]?Y;#,V=+
aa@_Q9Lf<?4BFBT?-feR?LTX]UWXV=3GDd5=?Ua_,[OT]M[P^JJA)U./aEWBGC>6
Q)SM)[D(cKCR<E7IJe#gUB&.4>Kg4Ab^IS_D(/cgcC^g4)S8QFg([Y&Og3M[C5#P
Q?>d)>>@I:7aF4Y<2eI><?(I13c)BR;JeME+SF]U5U0#W\>(&AJb]KHI[\\D2.<L
:bILeC(/\Z,d.JLXUO\ZECBD\<59WN(4#cK_R)f;L+V>59f&IUFPA)GfJ9FO;6L)
U_0c/@#FK#CR4Y6\3.)H@NZI,8Ea1/1D/(CC8W\.#V6]VgCI<E=7&D#/RLI(6LSB
ZM86MB@L-ffN/7<g-&ea84PLSQBbaJ--)A#3K4GL.+ZW5:HS,e;UG5I]NVf8_WcO
1?5H&_f2LHZ59)7)CMgFXJHFBP4fN46\NO.T;a&-+)cc>2P+cU#YdBbB=Ld_)-_3
f3#A&TG7W9E\;M7\W.+EB3&=<g].)Z)VY6)3[VdaO/bbNFJZD2+Q5b]R#2cF5V6K
C#+4GAQG:^4#fGO=eXd<fa\24Z1Q_LE[8]:<4C^,VXIZX)>I?CV#+/HfD2Y)>6Q]
M9G2^#Ng4IVC2f[>TCX)N+81e:2T0dgG/0;OV+PbZePO&P<_^HWX+(dQM7eV/FD9
b:fYFKB8OP5d=3-)B92AW@(SUc7FJ17Ub91_B(6Z>d,cZF-bCP@O;=Wfd>2YZ7C)
;2g+0;#?RS\UfK,R[De/GV?8<S7+D=+<]:7c4a6@8_UHbOcD6Zd(DF]5N1ESDe)a
_1I<aed+X6Vc,M/[&QeXf>@RSE[_YS1W[=0LQ)_5<PV<eRS)@SN20\PI/MfV^,+@
QD^E]Q.bCCd9]\Ia0?&YR6]&67ee6,1#a^#\#Y5HF8JIe[VQT^8MZ.@e&8CKI8:;
2PIDQ[LHe+(MfYU9&>+O__U9EfcQ-Q\Y4SZ91202G2KeAC<54Q(OT4@VJY^FM^]D
c-^7g]AR+_f153A&\L)e/F4PQ5VM3LM\IBXG4X:]BW?Ib))WGYaJS\37bXG4LM7M
T64W[#a4NF=9WV:8/XWYZ:ScY0EB&GcV+dT(<d+>f+\?4D<V>0=9/4\#LKO5:PR+
F:94302U_;8+DNUbP-91MO\=Z8.^,fB]T@Y>d_>//;fc6-5Z/6eQ?2^2>Y7F.Z4U
PRY@B9S[B;@Le+/8A1T>QQ-3I.d&:b^BRV__,[V<eR&Y;3-1U:eb3Xb#&=AKEZda
7R?LT@(XKYJ?C>Y8<a7-CQcfUYFdL.fbRE1Oe(65\:HAKUH5bQcAFLD/U,c@9USX
XaY#?F9O@gB]6B]G7Y&dQe(<>O05b0.D73YAE(UYDG-/XH]?_@,)P:4FF[Z6KV>,
4S[XId3bD<(VX?J-S#)@a71cZdg5dF;#1^8GfI&a.=+ZQ3),KW>2J2#\V\Y@=<Pc
72-Z<\CGO(XVOgGQe.eA-8eg0a29&TBgCdJg[_B7gb2X]aZ(<cZOAeeF7F6CfR,5
2cLPV&5Z5Tf_>B.H;<Aa&ZX0O-M1^1,P5-\2cO^=/C:2YGGK<:0\I4B^M[IX:IA0
VDD\gA3?XL8B<bW,=R1\G(<,I/W(+F0=?KD[g/N>LT?GaeJE?3#d]BK[_BKS]B/E
-#7PAgT;>R0KL624;a#L(B_9V__4K)/?:;X]NZ6KVcLgbZGBRF/C^?CT)&e+GA71
7GI^JH2==CEW<2[G_P/6,P4B=RI37,&7J,;VQ6.fcPRKaLaAC[,)LPEI4@f:D-JL
H8,.L0825:#D_Q5(?GX+=PPA8+>7IV-I8L:Y6ZYSOS(5;9NG^E:ca@1^N^<d.;<>
P(\KK?ALdR?&9Q1a&VfYOQR2Ea(>;9a&YaP76g@FK.:&O+\/C93D.PJM6MAOW/<1
>MR2@,G)(&7#0Z.gcU^Q3C)2=L?Y+c)6ZQTI<5OP&f+_L35E2GT(Ve0DG0[?[e<2
W+0.FH]45;-><YO\:15#\&CND^c4=?3O_@9[DZ=f9T:]8=6@AH7)P[/B6N849_)L
WdA?M&Y5ME_5I.E_KQ9Uf6W0MDH8[0,J:C1V/2C^adf(UN1eP_QKc<3]X>Ja(7<b
=WRc#<NYBdN2N_a?RE#,D[_SAF0gJ,NO:MbH=Ec0@c3PDRa\9W70>ec7\E<^N3DM
3da#5R+11g-<E,1ZG(\;M3EVD--^OSM8X9&e5)OgX00\4U_e7G5I<-FUMOZ#>T&7
X^8QFD1;^]84C#&>8Y7G\Hd<f<4HScbC8I>21G:3(I@@]7\=gQAN5=g6[43IP\?:
bWUW\[>D]WfKTJZ;d?YMR7,?+#,\2JGT/K=UaEUBIT&^FD[H+F=&b8[3J5B0f-TS
J&-EEB:N8cM>RNBFeVK]@T9C/U7-[LSF]<Y3Z\.5F7(Oa2ETQQR]8A/V\&dD;;Sc
>Z2P\S^gF^WA9H=7a>Dg8B+61AeT1OFV=LBTFA#1ZfSJMC359HCT(PeAH]<?(]^A
OdH1eY,b+GNbD[QG#,UE[N^HSK=V_F_BXf/.Z)dgE6bNbU9^1L=[7R\d3TLNWVX[
4c51V3<>7-W7g;8800^F/K#f2#13AX.084A6baDA&=]PA0FO;<,?F17F;T-U&0VK
^?.fO;e]0:0@+d/0JD>cCBJ<UY/S?S/Q50WT64fHP,eH5-2&>JW9:7+X^7JOF#5D
.CDG#:+]^VTLU<@-JH/8AFH3;7EU1eUX(#@BPJH<5g-0)1CMUGBf&RVaQJc04P?4
&STe^@1A+NUM27CU,4G+7)P0RM675gZgCORG&&dO?9O/J+#eUaTJ[O?3.:L&)TgD
.#]g8];W\2:.X(6G;ISZdC?;UV=[<]3C8V87-@Od/3Z#T1-YfF4g38-5G)M?:YYA
9b[[:KdHf^W&K.7AYAaaJP:OC]dZ3,2QH5Of^THH5R3MT,PO0;2<Y(>BgRX7K6.[
[cOY/bQW[@[XB4f&<9\YB.FZ+GL>[?YXZ,5<Sc^DHaTF/QO.:c2V4#MGC4.B#:CP
#bLEVTP0#J&B723Y=_]H2eYaMSD=d>E,cX1(>=Yg6Ke=7fIYUfCV5^V@,8X0OLXI
U5;G485SW#>F]&FJ?+e,ECW0:U3EeCA?LLXX[SfT,+LGD5Ca?+2Ig_#4g?<-aeX1
U)2L^OFM\#VFN(eF,&A9bX:RdE_K@C4H/2afEUX-3Hec2PNX\JISEVFDR?>\+_\2
C)bK?=P02d/3S<5?Yf&/BP0\&2CO?^f2d<7DK2LKG/CgWZ&cY<d]&V3/-b^cJVPU
^06MBf.dG@dE=>McA/4P^FLLH2&C8Ng1JQY?f(4)F[F^HO6G(EVAA28_31S.TSb7
?N<34W80T326-@1STeYJP_Q&IOCCYJU+gN(D&P=SN;>#f5HH0CNYHL?8?e<3;CI,
9\Q_dR7_#YX:#/LBeP-+TS+<NLY]48OOWPL9_R26DR9Z^95Gg>^:XO@2Z;fO7?]-
[CYX#XfLECPMH404aR6W()CC0>_d/UKQaQ>0I>X5S&dRIJYDPV>JN;.QKUA4U.OI
GH#2FBG1,&5?-/#\=W&&BZC5B0PXc2TD/Q?@Bc#c>f/8[MCa0SL+M9VZ/]/9^A4P
;/@\B>K@9]/ddR,Fe7M&)YFdIXX\-YY:\M/Zd\GH7+FTa@>.X(+Q?2Q=fFRPN7_P
M-98dQ-gJ1dZ=QKLHfG:I:,_D(LVfJU>?-TdU1,7_H]4V-Q)e7P0GKa#IbL@Q9f,
;+;+)cX)M+4aW-TSN+1HR=N/XM24H9;-df7Y3#fO6\SQcg6ISNdIZO;?1G9/GEQQ
85Ng62MgE^[bF?c:HD:e=@&+G]c@<F)g97S\d3dY&3EQ=4e1,W[RdZ+aG(Y>VQ7S
-<&:>KF0R7=N]SeE,<VH6:\;?7?(T33&3;,JMSJXfU@6ZX1.W;>B;Rb\F<d(?NNN
)G:/./+^:PG45DFE6YR2T=T1BOgG<D]aE9?+F\.2\P+MR-\+QN)a@&/8/c;>Z\&J
68c6/,g7PgXS:JSag[bU(HOKc?\,^9UfJ2)RNPg[--LK>2dGIWQ5b[&Gg7]CWa2#
-aUHC?9V?Z=XL)W_A5:T:-5Q>,;4GM(J6>X.&cS7RYIWY7b+=KWQ=OZ3U4@I1T9/
NI?PRYOQ\.8(5Tb^fJ4.A-]699Sa93^B9>1Nb?7A+U,=^0N2P6(_P>cN9\(T7,@)
=:2/=(2NC/bQ=Pd7<3YO5<&[=DK\RL2L8gQ/C,Q>Z4,JO5:JY]D;0&+)3/E<?YMH
SJ0]OL\<HN;U0#&B&N?N\G__+bJbRbE@Z_0<bU&UL:(.23LJCVa^?2_5222/AQgZ
87PJHa?1]6aD#[1&775V^17J=Ng^VZefd32eU4&bJCB7729^&dY):2+Ee:M+05eE
1D[IKRPA+]73?86_DV>38=,B(Y;_d&UTg@+&X_ZCCaN-([SL+2QWV7XOSY3b?ZPI
MY#)AB7O=1Y3V,26-/>\)66;JA.\,=9()9UEEIY84@U;:]:#+111_DYbfKE9OAY-
O:,(Z<QFE,H^:K)GAIeXGF:2a9ce>EFS)NJ1(8e7JO#5JNEeCOA/:FWGOU7gC,L9
aU8>.I:[LB;@CD7_N\df6&OM1@5^KG:[+7Ve5U&_>G<]^:D\XNQ\aUJR@(2;]R?T
QeOdNH@A,\@Ze0bK[1Y4\3GUFOP)3c1N?EaQ@VZW\__C9#3L;U/f-Sf9;18aLVD\
<84dI<MIUcVDg[?a8?BbfRbA7/G?)K?Pb.2>/IQ&+W6F,?fgM:_d60TB;G+-56M\
@@X19LNICV/cUBYXY=g5FC#Y(A@8;],N5?SRQf17WaYDABc)DMF#Q\bY]?c@BLRX
OadP(NdTEgE(IKPV&;W8M>>_:VL]/VV1UJ^VgdR33B<YXO?>+DXXg+RN1.-B7U>I
QF93:]@BWJ4X0,=MB[GLR.@1<4=G=aUU1RK5WHNfgCO\Vd6+I9-JND=FLD&bb&K/
N;C8Z/cGf8)1,f3)Rf.>cL1?7gTKK<),I/4TU#=]I?]Z>(5YQ[GXfg,-]>25=SV5
d#8-V_YOXa5)U??0M(R0\J^I,KJES>CJX3BF;YcQ[BBee&;bC[X1Oc=Vd^5S(LbY
d_U(O.>R,c^\[5X?(=51c(^Bf[5JXS;bP1?;8e\B\7e2C\YBYY_LY&QD.<6&OX[V
4@+D]7\A6LPe,F.,L3FcO83\@N.OaN=K?gY_<UgKQG_P_V:-NbUQ8XBIW3(GU&H8
MG0f)e8^RF5Q(:9?P<abM+8\>?1,E?COY10O^O.c^ZX:Cc:F2QHDR/7(_1Oa\10E
ga(M&-MA?dZ0g]=BPN#R([8&<T4J-:W0F>L23^/A&UJGX_7RB#aa6-KIF_KSGI(E
?RG2dDIK(Xb/?9=@JM5G?27P7F(IC@e&f.>-a^[4L3)aC1E=,-bO8>7A,gLHX2()
UdcHX^RAR<\>7aNL>ON7J7NR8<-I3e3^JgQR4,,=@[<.F]aAW^@P#U1V4Fc2/O+8
EcFF<?CT<I-0RJ]R-;Q;IEH6#JV70W-,+C2[:<@(=1,BEDa[BM^2-W(^JH2NZ9YU
DE]DefG3NgaG.dAe?)AKUI;J6@,,\WfJ8J5^bgEJM0C?ga9[IE8DEB/fd,+fHR)G
3A&<J1Ve6DRV#J5XGgQ=?LJ]2=JHFSH(a2I@TRJGc9-&L:I5QEGO#3Z5d6HfG#J6
0_/4SS?W:Q(+0K?P9e+F.VP.MUCIKBLNYgV2F80cb/W/I8:(K_;_8/ZVA;^d4.^b
bQXX<3Q8.a&eK?Be8ePVA>C34-(EcW2CY;:U2?;X-g:,.;HRe<2&?XP-O/c7-]2W
H+f888,AdRcF37aHR8_F9)4U_E33T44E[NF2A@8c&4e9^+&2bNeTYY^)SQ[38;4\
+;4TEX36:(N<R-16C]d#a8K_-Z(@^ES[<_@]J/(8EGQKO3S4XdBcaR#YUP^g,RbE
\+JPF1bKeR&H?H)Dg5&S0#<>U[#[LP]JVg,E&NG]I-<>2E:9?D(RNA-A<&8IUa(W
OQ\/2<?-F]G=fD^a]JX.fG/O=1-aT4JK-HSd>+RTdedA4EWU5QfNY6/D9AUcEASb
CC]=.Wg7>A\W;G:[5Z0I+>W)GDIB7407AL_eT]2ACN4g[OAaPK,1O:(Z.Ka5C]Y2
A#XW9DEL^R6>O(B/C(:;.7P1&HN[aOHX]eB;b/,KQK0d_+?GAQFA0&-@L?O#QVR5
_<?];G5(SRZ&YI9Jg#\S]0AKJ([bF@#0?56Bc-2PKYc)FdO.#0M-0WXHR1]79,TB
+IAK.\ffYbHUV[[4>_MIA&CgNC&):\YCc]G>bR:D+JW-+2=(6a34fD9A=7<@1:>R
)-cW\&9fa\Ee(b@S:IJU;.CA6;U5,C@DY=fe[:cYGYf\aUfY>^b=A;c5decXJ343
9O4AC:GW1)VQD:W68GU,Ic8M+T<V.^<H^S(gcEfM1HJKTdTXMa\?;a/\E7C(:dMP
VO1?<FKf7=PA-[0/Oa44R^BV31<67E<]Z0.e0M>-QbL-&PZPK)?:5</N@1DRaP,-
[R():C2-eNK,_H,_)2^+P]@84S._:/RCD_/TL0J3.L0?VaPc?]=d9ZWDe4J0U-24
7[I&J(c=eZ5(R[K<b_ICXbVF,DKBHPY+1)Mbc>aN1ReK(<Z370Mfd^VV4T1U<\9g
2O9D>T]G]<PV)V0/.YeceUQJ#P\4S,_OKSZ&8F:O:_UX=]fI\Aae;IT1LLON@U67
H#5]C-/cNQUR6J>T/:ZaQbA=YC;;5:MG\[/:S5f;U,.78Q,?TcQ2PTIP4(5BC(Sc
)K0Y=T)XRcbTMYc[V4RF,9POGf45B0<Y7;.CPfI8W)+/7OK>])_UTd]NOR)L0-XK
+UGB30@5ge;8@GS9J][O4@ag8>;4,VGM6O5Dd)JP&/5+Q)aBG0CSS<@.d@ORdD#P
R2_DF;WD]9([dH1BM[AD-/AT-(FBWDEPR6<8YG_CIbC>=YbUb#;/bD>.+7T3K\M(
TK:V]OEDZ87KRS3K[:AZL&DH)XVB:Vb86^MY.0MBL<0g3T7,#7A/6T:&Q?=-9C_+
<&C6+L[7XO/G8M+H,;V23LZVCY_gHL\a+AX@GH31MJ<R8PdE\^Rf96O?DcX=JPH@
I;313#<LFB)a/^QL5[1+#dXL:aDf=@O,C1>(c7Q(W9_:=;5<LZ0[;++.QAA-@D=F
LN0[+04gS<K]_H)<F3WAA+f>bgg8]]R)O<<7,MO;5OY^ST]ZgD)?V/.(0_[F</^a
JIg+]S7>aN@e@aT,WD#,7DLc4T120-RE\P0IU:1_]/6^4?_@U[SC]F(1K&3XQJ6-
R2aI#FD]<1+b.#>;<_)WLUMT]()egIU\)aKT(#U3L^#TbXVQ=;:(N_cY3aF2MgZ[
D1P5G_IRKBOH>B]AO:Fc^#W)_eV]</?e+Sd&J0Wa,2:;WR8#&+ZZ.eG\e>E^6/AG
Uf;?J1P]LXSWeFQ\GbDJEaX>9-?9ZfED@]&)3NZ+<9U8JX?VG#)?Y_M7,QCO+PS_
dd=TG=D=aY\(U_>IX^Y6#/1^NGbK5\_S9JSKJ4IM=K;_)eP;51c1.H8FQ;RUC=0N
M_dXfPa\<QB_(7&&PM_)_.g+]6K+6S,FGPGZ-FSFV_bbL/:QNRJ+\MNLG57A8XY#
#W5QeSNM[Af88GI>CRbV4c0PGaFe6@[<2I=CUA.a]d&V<R;8[e=Q+P]5B-\bd0,L
;>]e2C1g(2-3&C.f<<ZT2G>V,UE-CQUEa;^(>W[cJH3e;L_B9UR/b3W/DL2[ILG0
ANLgX/=d4JgLZW]73T@_&C-DD/.S(C-=YRaJ:,F7A^;GE\aZ-:-M@^,<B\O:Za/9
XF:<-)e(=L_()7U8/6?C>8DV]fV^,I5K[&+W1,=+e#dV<J[OIM7f6L0AN-Z21/dE
JfGPO^f\W1a]Vd_XA&c]\e.BAg4b33P3&(@;FfDJ:--^a(Z^WB6@5X@>PTC<A\5,
J6Jd<P.#Hg0#.3<TFP@[DJ]N,W\e)PRX2O)]A)NQOSaaZ7J=2.8/T^LdTgY6#a(0
-c)eFe+eZW\M6Xa>WgY?SHQI:@5RP/-TM.F/].BMHL680D?,BU4d4-H:4fE<#LE(
,BC8J0.]S26>V8^_=LD_,2PZg40@US)GdVePNILC<71VP#NaMR2U&#8]d,0FZIc<
H2cfX#?gg>VYB]gM]S3)8HCOKbe-dN+?H#(G#4P&KSg-<9#BK)Q0DT,9^6+a)RF8
(5-,DO=QM60+g3G;I1FLI<AQ0)\=1..P]E2^-H1#:-51K\M:A1-[B324^5EAECF6
f5LT5A=gDST=9G587)eQG@+JJ7+#bBXddd,fTZ6NP]?8M#cK>LWCNL_eUT1NRRHa
L4;36(F7WfW@RA][4f5GE.[+0K_Ze:Md)f@<DDB=Ye)RWS)c9N&0U;L0O6O[eY0<
Y<(B2@XKfD.82HY@N@BV1&02R<DWB?T])@?C@2;3LU,@_^Wg^W6=10^+FND?>Y/2
/B6+X9#O:dI:-NUXa_H^5#SIB9E03UbMOaTL4@8VS17^=1_<0VZDd.H?;4YJ,3+e
;-1DbXG?,ZAML-,fL8JGFTaU]58^6^0^/)dQ;\Q9SXBIE2994V7#8K30:T6a^3MW
e<)-)W:RQ\NL1fB/?/0]D1^].L)]/RX9XQI/ebgaAFKU1PB]ISSY_eGG[N_10e?Q
BR-4E3#_>Rf:g6Og3BQegGN)D;eYCBT9gc_@IHPVX=>aXV-f6VD?2DD,URb>&]1f
c&4WdTaWHP07XEDe5)4KEGE.>&<bSXR3Y-Ma^I.M[0MRT2BfSa\1(=A3a0DJ9-)Y
.N^\\=RGV#ZRdC_,AI?O:P,PU?bC4&]/CBAW?>Y0YR9#=P1S9[,1Ac)E.8SYE1TO
/#OWZT=agb>[1V5<&U:)BCEb/+WCZ6]DQA9=8^./a;U218&\>G63#IFNL7G/+<,W
0C<.7(D-UWS\0?-5,B\#c16<c,>M^]71C[6S:1)HcQ;3@APSd@F)Q;SY_=U[)W4^
;]aQ58\V>&E.MA(Hd>X\(I^c64f[<c&4#,Ag.K@-_bI)E/U-IK2V^=VKdJL4(-Ne
OdH1X^EA:e>X.7G7K#Of6+1g_9@M#QQ,DbW5@eeM<:^#b#We(G7Y)Q_/>:50;4=-
FD2(J[6Z(F]&2L[>]42eIL@F9a3+R<HUfcJVRC]GePPBK9[Dg^g3,B=N)@..Q,UM
[^@AcaZ--SS#ZUM-J^KZe<EGNQNWfIC9NP=\37Y6:O@ZNV_gR#,0?S@TE\GgbU5]
ZDa]U;fIC_@R6XgP]GOLa,U-K3\QE5,J&01;.B6O/->IWAT3Fa(d_M4/R&I,\T4<
WXGETQ<F.D\L#(A@K.+Uc80Z]fU;V?;2>YYV&MW</^2Yb#]U85BW(T\<N;5e6KWa
AD-bKA7(+N0]IW?-H7X9#Z-ea58UKf.Se+ARaE^MSA;IIbFCPB#MFXaQI#DJfL9(
Ob=T?Q[H792-9^A6^NI_C7N--+Sd0QSWR0,)Kb?FVZaN.#.ARa_]LP7)<353D_@F
B0/-gG9K_;S^JF=W5Ea65&RO?FDQ67-6X4.-eQaC[B\<:5XfFf-52@;YHSR-5SJ?
O.QX5AOP8:A>3N.R@K-3K[Qf=T[#/Q]0FTG-_2_1,#.5\5+VG\9fA^>5QA519(X9
^10W+BWVFTH3O)3-3C\3/&WcAKQX61[,MV/01RA[4g]BK3E:8+fC+Fa)WA[FY;1.
ASP(9)<AB(8[ACI()0,O,;IZ7[M<BF\W>,JRO]aCOX^-HbNCdS@9/S#8E.XG5BJK
[=RD;,KJIZDG+NQ=U)M3TMf^HCJe\b7AWJJG-/VXD.&AZD0d:NAC+M>_(FBX:#N_
bG?920;9JAWM+MT)/N7TGLMgUeD48K62F6BadL<J[W?)d1MCcHX3TXb/7Q?6M91>
/4HMZJCJKgW(VLc#3CgM(^e#^M:(KC#X<RAc1RI@TRO9N#:/DgcEE(OgFNI/Hc>I
28<9GUSI+6K;[^=:KS>G)#-a9,82P,XURG(DN\8]#\::KG_Ud6P?SPbG317YX:S&
(Xc5[/^R_[SeZ3b(GL9Q.J&V\CS4=R\Ae\J#MbF:a6:gKSZRb0KM_LVWUS6\bQ68
QHC6,CUO6e+Z)fB/@FBYaX?.D<XONC0^fI[@ZT^Xd#E?^KGHRB6O/Z/F-.946&C&
:F4UX55YZN?03-8GUL6aR+E\:CS4;T)FP1/.I#]BB7g+3V.RD_=BMBb7-Fa&/32c
(6L,LGFP1NR^7&?V)[L0C)N:ZI1@g)d0eP@Q;PP9ACJ;6<&[ZgJ24SCDNUNH:WJ,
<O/O;YU7=)8.9XPCU/XT=Mc<<BN5IV?[H3ed=JAY8g3(7&H573I\,Jd:<U+f?/0H
HMBf,8+D4W]:S?I;<Qc2O6g7EfE&>dGKaRcWPV2R4Oc>BN-dVK8gc>UC^(T41g,+
bIGD@T#GbUd(Pe\b7/a_K9ZUW,Q1CbTc8UA?PL(V+_3I>M17XT[T+L=WN]KFK^XV
U\T6X(I>#0>R3_SJOY26PdZfGJ=?_ge<U&RgXFc?+HEHU>G;:@LJ6X:g5aNg@1JG
YYI\#<&0WSPHYP/ZYODF81X7S7E?@GUT.T3-^.+D(38]-2?+#S(>f<JF,\[=UIdc
]&+A&?c]/?(YIXKL5MK9>g\OZU66PdC<Q?:@cg69L94D/a-FCLg[V9-#ZJ(.9>29
9O9cHI;=Z:3)ZSAVXZ/.RBBPb20L9B\01&Fdg&]3NbE)UZ/Ig1Vf^)\M@R7JJ/7b
I>)1+P1&ePL>-K\X?>5>5598Wb8#fYaKDPXNLF^Z5d[XBNBMPXUZ-2MCQZL&8\1W
PE/a1?bEK<)e-V.JC2/6IASOYKCg]+SbZ7M75-ce:fI@I;2I8)BS.HR9?dXU(Aca
.UI;35,]&B^(X;9<R5XLR\GM]#//2M[CM.65G\b6/(NTa1bFd2M\ZYY)KAcCGe]K
;&^AEEc.:a:8;M9U@ULL9LIWD,\P[D[+Sc9)<N;//Q6dS#3:e\]4-0(@E]I&L;-A
VFa1dO;+BZ1AUEXgB_<Z[g5L]);g_P/5e>8(#&66_NU[;R/IeI,RUI2I7Y9=SE:H
/[VgbdfHNH/.<e#CVR,UL.Y2:c)^/Cf4<4>abI^ZFRA9,>B>=@E2Vd[DB>;</g&X
P7,7DN[;WRg<=[.S\QSLdEHR+]4Y&UP<DB29UbGQCS/G;b_(6ZCJH+B@IB9[\&?D
.3P<96__Tg7P2XAKIP5I)Y_]1[e4V\9UZ(IaYF@7ZgV2cgTNL-G&=E[+ggK<XKEQ
&?,KPD:[2<Yf_>[COOCVT>>^QTKY?/73O6^B_(UVN((?N+F)5+[LN<CWD(Xa;6-A
28B);N7=QPV8WQ&S>(I<JC[-<?]3_OO:.)W,F.6:Yd4>YIEH3K&=F-H>]B2OW1EJ
?fc4<8IUMfRB\//+E)0)W8#P>0R&0WH.dJ9[)GEeUC\/IAHL[T3#B:E_Bf<(J[La
B.Q?E=(b&S&fI0FE]:71EWYKU][f^3OTGA\V[G<>=4dC.3EY+5K:g4-<^gC:673,
<[b5EA4>=D2?R[+UAWK&D)<)dKJUXD?^7>[aK^;@@+4(CVN8]2IafZfJ3Ug+HU-&
:e0G_C0Md4&eAbg-e[Sg&QcP7>6C5NWPKL_U@Q9IE:cM:YKMZH70NUZ5K+HT8,M?
W7:6=QP1B_6bZA9BA9bU06KeKN2N>S3I,&&[#R,(fM[EEYQa?TXA>c<[UBO)Xcf=
Ae]f-dY,_S-E[0;UHRHO431/G<\E2[C<SF5X7>/6?;8@WWPedfX7E>Q/L[]#,\JT
WC^eA2fC/Jf2R<]OT=@)./Y1,48eHa:&&P;)3b8WJA]6fT([),:fUT.PQ5W6]EA&
a<fX0W3XSfa5N-^Bd:/U5-KF),YD][?(0;]g<N?^G_+@_gY4QN[fPgWM2dGQ@+[>
ZXP[)>MS=<2?L/^MZ2\W:@Ja,Ye>Y2<baSJgIU[7be4dVXK8?f0,C6gJBRTOgAC=
8-FY&,c+.MHHK-UBO:U1O3dIM2a=EeHTLg4>88)OfY<1KV&RGWVKbQKE^ZX?)<#U
^Q=g<.=X>Y<<S=<LYW#=[g+g5E4,8<eW9^\fLg#F&dUX5.cYa3]X?35e/?fMZB4)
&]3bXB\F;JWF(_/\@YX)#TL5@7.3OIIX9X]EEWDJ9<=;>ZY2Xf,)=8Jd46fLJQLO
^_=6I7SgO3Q)DG_/6=&T1<1GdVM?V^@-/1)7.Cd2=A:23&J0:8PK2@J?U)2ZH^>M
Lb2cG+e99DH4N]U>f)]Ic<cT#@c\LaC+Q\Jd6LQgE=R,HWQ]>P246NbX7H-7Ye7f
ZTfA^&-.M5CF;X_M(]S3O)3dfN)70>#7dAY2QC.(]c@b>P#=^0CM/f-6=5@SN[AZ
<bLMDE:W4BHQOY7HY;GQL_A8JJb.-/]/Dcg+8Z?bZX?1LIIfJ+S6[[&D)#+O7fa8
dOgEQ[1cX??<JX[,DXGSLKaJK<+:]4JgTG=Cc0OLD<.(AM]LWc?\)M>YE,9A6^C0
,(X@++LS6Y\c4d=aJ++1Oa28[+PS_U\2&A,:[3b2?N[\;eRCH@b\1>7FOTaI7O/)
LbDIG(3MJ=6ceP?e/Q.3CGD7,#9EET-g\+-7NIA_^dgT65[DHB6MTR;(+YPQ(=cX
0,)eJV_J(Y)^HIQ(b/\Z0Z2XVF-UfRA,=@&g4-8\bgA1KRbaYXNc.+\Ab?,A7C#4
OEeP)\<g1JUN?K=Ig\b<#?3dUW<040aJWLOe6]?IaUW5JUHI=]?>+>#eSI#17Y_\
,d>]U5E+LMA=]AcW&5D48:-Q1]]gaCM:N^fI?1/+K4\MPS]/G6K7I[f/cfLU-0DT
J&NZgHgY0\DLd&c\4S_ZfXTbf=U0N+:69(\13&:=f\aZ=7\+NWMK#0eGYR@]_[AL
^-@<:BBN);JeW0Mc2W314;WfDJb7XC7/,V@&6\^92OZ<(JQD):eeS5fPD_O:/+bf
V9AK60-RR8OY)_6#[+4I@<HI+33d7@6LG8<^<:(L^bK?0CbE#+LU]bU45+FOI.&&
)]F6>DQZ-B+1Q4A(M,eS-;F8eNLPO_^ZMeSTPFJ/#b]/)3X-OF1G7P^CbX+?M_)2
ADfQ<_C2d72.L57JG0E6)@D[FCRE;eC+W6:W/?9fLAB371,NcR^F@&8cFg,#@b#C
)VNfVV=a\D_QX:51E_K<KB7;SeE+#;)g4DbXUEE#fM:SAAd:RBU8Q#:g1ER8TT\R
C0c)d:+TW3=+aZX[6fW6?1-QQc76B[+EVJZSa_f?2bP6N]V]+YHGA(]82EB<0b,H
D^.gWE9[+:.?9)CK6X#V<MX2)bX\/C?5->f^fMGQPGDDL[U=KMQ@.VR2d(JZ:\:W
(ZS/(62(Y1C0XG2e@;DYKC^9b8V;[^4,JT.?LZ(5/6Gf.T^TI82\0ZU/)]7,W:?0
<C]TO9)JOTQFd69FZd1B+=ZX^L-&O[NbX7O;><36?,,=Ga_)RMPfTB6b3A.9c5P;
<c1W,a1O-_/eIgU#cDL94L#4_gae>=JV1Q(10.gE927LD4J.I]b^VCD?I.;&HM-H
4dOVM,[U+J[Ua28DN(MXKX=]_d9LMTFVWe[]bC96;:#6Q75-APWL:QY&.D;W9U9X
a6+?)XDK6QabBc[.(I55b1?UD1S53>1UI&J-C@0+SZ\)>JL]:<4=<4C]UQBNFS75
PQg_DTKX/^C&:d@7b=ULQ\g#0_WcWJ80f+_\U[7CNLGR+2b3^=[\WH8DXbY8f].3
3If[#ZB-H3YeIIUFP?PPH(+bOH27=WcDO-?TQV;?F920@a#8R2X-LE7,dbY)8?NH
Ma73fJ<D&1ANUVGT7IdAJMA<32LbfeI11b=-3bY^d7>]PFJM>/FaJR36:]a1#d9R
Wa+b@d_]J.^=A&>Kbe/.VC_O)1,8POG6e2KZ=;,UJO09L@#\U\AFS8PeP/P?>IKA
<-A\Y31:FI8F\LaTH)e&#_:d,AX44Df&6JVYIP85)?7:C;WP^NY6;0H2d8J+5A7P
JV&+/)eL]7V0K;9IK(>:#14g2D-^Q1dKQ]@S,f>3;=:@T?QNSSXC^cg,H)BG_TF?
V7H/G]V9#DMSW+H.2CUKRYSbUFBY=LRLcGdY-YGZWO=BA.T@>00DYe4C1J=T@g0T
ZT\eFZ14K582ReZV>Fe7bQB.4aHED1:V6L<B+@9TFFJX<1[R[F;.^6^F?4ML7&c#
NM5ca>AcX4OUZ\+XW]1/8NLGIOAF/@8b94ZN@cV@2)5?H31dHUPd9WYB,ZKPM+>X
d6[R_eE]0/^:WV<C?OI-<36_b;G/FFaQ=CWeLNNB3Hc],Y]9LIZ_-(&M/(NKAZI\
4,KZf8:0=]C0HJ=0e]Kc9NZ,ePaZB=ROKB;QO8QN<5fUI1QJA^M:Z&Ccd#EIaM^N
RY=RN<XfHP_?gJ]We0c(d8UTP]X#.]S>&M=/DVfC^KTQ;eK.Z7bWK1+O0eTcd#T#
[BC-Ha.7VbD)TIPXG8V/=g+Cf3F1#\DaRL)N^:BYP+8(.JQ\5H<(1&:\A:,>BO)T
9/<HUW8P>2(Cd9Q37@B6c5&/9>YCc3b^ON#59P>AASC)ZZ?A-YGFE_V1C.1X@^C=
a>-\9U=:965/@;\F@gUE1K=_e<(LE,e0(PVR[T?,]QYD.B4]KX+9[\3dL,?&L4ID
(A=,.A^WLY7;B\^1geJ^]P+f-fd^.E<[&,]LE#5CXPaA6.bSe4ZNPHK1JN&4F&X?
#J?YD.NC81KQCOS7BP@eW7RZdGIVUeA:D7DFIW3V(:TA1;1eRa,V)cd@HE3?BMW:
==E?99;GI-1,)>LO8&S>-BP-B<;6+=gNYO&fQ<WL_b#CU&-PcOF+MH>aVS_0(a+K
d#Y:[QW=AS7K>WIMGX/543K(IS_O2/_bW-^@f9(&dI#Ibg\>J<MabI-6)KG@9+47
B=?,GC1))N0@V3N8)P@E&VNW(,,dE1d4?6c.V4^d^^=NBUWU2]9TMX9:7U(=CG&X
+B]:X^3BU&;V^+7(YW+c].G)B2[UTK>VVDK?e;/PFE(V2C8;Q[9E(PZA\PN](<KX
ZUOLB98[&.;3#9LJPSZBZ;dcQ/C=Q0DTB?f(f&Nd[OEa)XDIQJ13GO/g&_JA1fFY
f9YUDM0d^TBIGQ][2HLRa?/1VE2(7[/KH\dJ3X7\4PPD0U,F+_.T@gY#:,9O/9,>
Ba4(C:D9B?/43H:0.Q<PcBEgQ&D7I8aTS=)0CGHO@.8VbK[]QKd,]Jc6g/.2-AU:
bE.;/IPbIGJ1(I;d_ODfaU4[Va&E&bQMNI:P)QDUF+JZ3;M.1Uf;K6;7+6]HP46J
9a=<#LD;@MC^:MM\e\C5KEA9.aW)EF8+]M1_cEKOd_7gdYNN;-_F4b2B?FF/U9KQ
c&@0LLdK;\7OB.]1Y0Gg^VWP9F0PSeRN;HO??+^U/aH@+71d^@66fe-E<:9cOT\S
cQW:\.g:SD]&?)4+3gRPRXD4/1fW5CAaV2I+=a5dOGX;LGYKO&7R/6V327XF6DJ)
TcR4U\\acfbbQ6DZ8N5460O2D\0([Jc/GXEIHWN)T<b)R#]A<H_8cTfX7[;e[cR/
Y<PZYX[d9ba<aH,eSe1H0=Z:W;U1JX,PbV9XL14W^.DAGBHeK7)ZF.5V4)?b)NE9
]1NG?&@(@e&X_f:Z()?ATb#]CCdD?I&MQB@8:Z@C.W0(TN/7B,)dZ@&?C>FIKE[A
4PYV5-g9CD@H0Ud2,<:);FLGfX&Q(0/gFCM@K+F,;81Z6d/PVGG.Tb8K0bZ8@5gV
ScRH[Q+=L\B,=87fX00?I_((Y&ed5MQ5V<Ze?+HV#MO^)UXBV)H&-K/4I\V2-B^<
KC4c=4[^Ae#a9^&V?_fIP#B0(2>?Q_cE.O:\I+YYaMd6(V(O0BBM,Zd=?E/=O\+0
V&g(QTU.[+4U5^HJZUC-)35729-)>[Y<RC70(>-+G-3MfAF5DT,0bK9g01R_<[<6
X/SMKL+IYcF7F3OP3:H+IT/#B]/=SDBdWN>VR[bbHX=L5&#/0:e[R(+X//g.KYL:
:NXM4F3>da+cL+[<;^<212-&&U&G5]b1<<;V-VIJ7ZIV;##TG7bE]F])VK@S7KTQ
8gCF;ECf[\.=Q[=+UD5J[S@HZ9LH;QMTL]28DeKI?1T&-&T\(&@,1V\1+6Sf<(_g
b+TUcGQ0OR?\:-0^(59X.OeXT(&_0QY5EX4b9@:(7Qg698>X)C)&B.#@OD/0f.<:
N<XHQGZ;?E5FUf7U_Re7J_<F7d0;Z;gC?=fV8KbN4-.dd^Z8?[Z\0ILGOOX4UZ[(
9EKXW5C4Y:bc,Z?Hg@6IM87YS4//L+2#632<2RMWS)/#d)g]G[<^5>T>QgVHW>G9
cRY.32UA95[g/,H7f\[)8-LWcJ&5&V-L#;EQ_LKf?.FI@^/=UVX3WCWcg=g;b[-c
c6(1<B[;D7^#0?MA+..8R_1,_-)@XJ.,T\;W]5cLK]7,+<#DME@J<\[8V2J]W+<Q
Fc:dT[LAKcYU/KVJCIc2UW#3&0+gS#Ye9,(VM<6]..;9OWGOfRFQQ>HP??C7eeWV
Cg<RW&QbgKLP7OE28+=.\UB+2;5dNH=7RK6L+DJA-<E7V=8\G2b_0&4-6,U]O=W;
CM8e^D9CX42OQ0Z<NcNOU^.\cNKPKJ>ZHXbKXY>KZ/E;VCJDQOgbQH]=4g<,Ub,=
TC9[UFc2bMO_00Mb=NGD0X)3FD]cfQAf6#9T\M1.>GKM_ALH?MSC>ff^-PGTA0WE
:H/YJ;;H<I[\I3]Kc#_@eb@.D#dJK-9fP2B]DgN9C@.C.ORZFH8(a?@c7dF1QGTG
>^QfaPZ[cZ,Y7GE[#@+MTO;ZF/Ja/FT,f\R;^+^Y7K&]T?EMTXf7g1+2dHL\6J>R
gK0)aT82eP9;F1OHWM;IBKb(S^.UK0:gW-eN?cEIg>K45[:[XVNK[3PWZX(gGK\T
-R<WWBO;7+J[1U7@B1HSdZ^6L;=73G@4.5<NFe6CS=91X@2SeT/\5J>-:[EWARGA
F.gB)BM2L@R_.A)ZR^+1[.a:F#XE4:AGW9G9]G^MWW)::&Z17_Yd+:VWP(e<cF1[
6>=AK,WD968H#U)HH7R)R1XR7\.JUL&<&\b,0R1Y?UP>>X_0,?;(]WPZE^4T7O]-
R9>@-VP6:N/)2;A@K4>++1f^4bKe3Y@(:RKP&OA30X^cS\VN+A)2(?.J2-U]Vf&K
[9,GA-DF=>^X5_U9C83ERGC)3=#UHU,7T@IK9-a_[P_1a^3fbO?-P3bB9&9.?F_&
6<.=T2#C&H^c^FUE@T?[YG,[FLb^&C7JE+6OLUOcARK3,(,G_&c:U2X^O.G49PQa
K)V.:dJg&CIWG\af_)WVDGEJaeI:C\FSNTa^<PK4XHI[HL)YFbH^\YgP5@&=+YQ6
DZ\DC,Zd&VS_eQ4:<Zc<&9bPJ3Xf86UXd>ZC27VR>@@&Bf?/IYJ5?&FDXY<+2<KB
K/U:L:T\c;bbO:KK0WdI_/J@BSN>>[gKK3,Me.OP#:CH[6MU<5D39H?233eeP<53
/;+K:9U_2e\#VYbLgbg@Ae@Z^LFW;\3?/^57K3d7UTDIffNZG@1].5F2bHCUCfEK
&N]1Q0KT_E^.I4U=.0g-A_9;fc868YSA1VV)S8IgLMeV+XVO_P#cgA+g?H&Ue9Y[
\>AT^0(U2]K>:7JAbYXAb:OO(5:cSPL9HD3LN[3.7TFO^)MB-TGV58?965?E5_)\
5EL)50]0>=gDa9cf3SX7&B0/)O+,S0U.=3?R&V3<GcT4TJC4]>;@Ib9OC/_4TKAQ
ag#a\E]g&dMLG^Y>8:RU2_NU^4U<6U(#8D\c7?80GEBJ8.T0ZY#S98LN@ffO?FSH
?H_>cHKII1X60Z.78H/(R5S3<;)D,HYU.RS&DMgJN_&PT#7)1:N#@a+<0RcRFWaB
cVYg4PS3><+3C-F^)bUMO#DQ-:VI^B(Q/H28C;S-f_1KLJMEC8T9N,b+JE6Vd\>^
,K4TbU#<9be4]aEgfVL6=bcR:[WCcKNg:4Q6F:O54L(XM[Y?6NT5.>&=O:4&DT8T
4G4cBb\fFYT0^66N2/f/EK9,_5;A8b,>HR+e_R0@#<)JDfM0Y:)V#^CNM1I_)VMd
C;5:MaTMBCA54>V[5=F+db\98=@WFI>1\=Y@I&IF+?IR6)b..d1&7K1-?f:AY7/.
&5CJN\XQZOW02380NfK]/9;ARC,JCTA?c,9QPS@;^VGfeDR9YJe\72_9K6JY,NY6
eJP0e+.OP6b78,)HP\8T;+[86&18)bPG)2gc2MA-+)BC8P>QB#Y8?Ig=&S\=9NbC
EEN5IbeLdA;b\S[(UN4>E>b[7UIWHaa9WN+TSGM2,^SPSS[9MM.P-:-]13+762aJ
4OYa>+H@\0<Q+=@->:c4^M_S4IF)f],FLfEWIQR(697GF8E@2)I,PPEHYF>]cBAI
UEOd)MP_aQ7SJJDLcBOR35\7<;OY2_?_8K(LIKU&g0Y2[7EP_JBZRYR\(#C=5@.@
SS.GU(gQL(NHe;L^5NUPA/fg62Z(;?:AAJT.[CSQD[7T()=L.<0G38+:##)=5=ZD
Q;5@S;EbaFYY_8UWd&)^0-OGFO/FK>N^2a8EC;9<IPG::<(DKO\]18+5:.56;c&L
3KAWPd?>78:/?G1#-K\8];JAeX(:4ded2?(QZ^F^bUK[^C(b6/9F#VNO?ON&4IV5
RG?]PI^:IaHc)NHV3ORI4H#YF.3&eM,=a9;VHDe_4C302RGS(_^:@FVJ.3#f/4P(
We.J37VWYTMe,,8=N5FO+^9QK4:9B>cTa3@^__[(cFVc=N+>L>/4@.d#G@[e=9-_
&.8+LD85b._8=,L015W[eY79gJ@T/d;7RWg4L[I<SfRU.R[8HV9@\6R36<25_d/W
7M_@2TP+fb9WO3fg\#7gM1VGG(AgL+\/3Lg#IePPRd+ZMLeebSSef-K2[c_AGW^S
cc=[.?;aX0eQCa60UW5CLa.NIf2.0VaXC03--Y5H8&^63c9[&A@_W;5FM_D5K4H^
[\C<4JS^=:][MES;d31MXAd]?<HX/2A<PTC0C<FeLT6e([,6QM(gdeaP>49<?Lf6
T>P1^##@\@=_YVDUW=HOKQ4_6C#RTd;#(b\2f2_DLHDZK@D-ae,\5IC@5UPdA2B+
d22c+M1TZBF186W59O^UMEeT6>>gNG4OCf1&6\@^\3\2>2AOMCUJCe:];Q#8,R?d
\:SA=dK/79;0XFY1[XTRQY#<,H[HLWG(R[.TdK<\V[\\Mf0IcJNI1.RWPLXM73(U
_cJ@4)/#QA9]3Bd/cS=[WKdDbM_&ILAQ#;VSOO=(K/XV,LVD2UNAFa.NN?DTXd0:
=f8U?R.XbR7f@FLf:1?/T9gV\,1RT?C3[MdL_]9<<72+dVEX:#KEHEP6DSK3I]R:
6[AA>3a4..2TSWMcAEEVRTD6[27BfHT14e>PYg5>>+#K+?,dd)]5#Z22,A7eaFY4
Q?^aQDR9H@XcRU:Bf[G/:VB-^TB?M7D(0>Y4?=3d6b?EGE3UQ&C#/Cg0c;C4].F&
20CONgRK]^Ka#<1KSALIWQGGNZ]3+d)Ug;;gK#C.V9,BQ]/9>ePHQKR=c=J/9SPH
H_d\RH?b?0408U=G\fEXSUG1[#fP?^?\NFJI:V@?)E8<<.7_-)J(BXC6.aP(Y7fB
U1c8ZQ)b>;1O<OA;G+dZ;e9#)e<@Q_P[FEAB(R)^=.JPCf]H_a2(;JV7a8=[e<T9
ZK(3<a8IeTEaT5[FP_e]MfNY+-dM?TDOR][/GE4_=<JA.cg,<ac@SR@c9_L>5;]6
dW\ISdRJ49#G[A.FOJVWZa/[.]ASH&TS@0fVTW:;AcX)>Rg7#76)3:HON2g?;DaU
Z7C>&8ZCR\DW4S#/g/:2ff<@HBBTW=DW,D\#CTS(E6_OCQc[)Rb2?67BH-:8W:/]
E4+-O\F;e-1&+Q>,XQQ\/UbE63NfCg,FFA1VaXZW?7:BU.BDg1[D]]aY2/e3>DBY
:2K9GI88JUN/<0K4I+3?Q4/K2ac?b/B&=MHf=fH+7,D&DRKR9LAW[&O>;S5V6dc.
c54OaS;WA4U1d<-]1=T\ZJBYeQY/LJ@&aN?T>e>/EE+b,_7_(4W9XZ-C]=HEZ^^)
HR6_A[&L51P:[EB_VBdM>^K92c,b1[=Y69GF@M\E)L_,7:Q.YHc]U.2Q7<][La7K
FR9f76ObAAVH_PAeJe5DT[C88MD,M29M4N)g3:GN&]]1D:2_E<JP;.O>bb]XYc5#
B1b-Q^FUG:Bdb0YX(\bIf(LYeWb10BM^abO,BdV2?2(H<e4L_L#A?X+Qd@&YS4IR
,g;G2S]REJZ68X,B9:0D/RE)C?ZF6SCG2+[)#a4KFd98GY^UO,G.AECR(#]fY@NJ
87HP7b:dPLd>?E&WJfe5:RBWNHH7;XL(Q7H2(J.DgWD5.JN5<M,X^,NHfBUf8&I6
=04.[/FFXR-3/4TX.7<46AS6=\(;EEHPLI^FH:Id7]V2Z<^6T;IVI[)6J.V7cKd4
G)3fHU-f@B>_+cg2:d6MJ>TcAJ_UDHLE9S0=T/A-MT^?bS:G^@TPQP\=d2ATUPEE
aYF;a:NHO:\1B.NZNZ#<FQ_K_5f8T]bU[8^V-RZ\CG;=&Q;WAJaT,9fW,ZZYOHY\
:^[Q:/AB:_:T\MR+[7=>P^+;+231\VLd5)MN+VeX]a-;7AVJOd@HNb[>#.W;I+SD
B0_3c<b#)\/CDgWFX01NFVf?D8_0=EJ<E]0W;GM,PKYQYMA(0\1CV&DL<0?DWBRQ
P0[D+J109ASBG[CG6FK]C,#^?+DI.UKaL&VdEFLR^.LC=-RHd(3OY<XQS<,V.ND^
Y@Q>9A(R9.J;/B4dK>ffIT>dPQ_0C9C]J<bO1:J+0@ZN_=5(:=eaAV]Q:Ed)C[4;
U0Q:<:cYfcM(D;2/0MKYDW-_TY66a3V#8#72,7=&29K#N8fI#,GI^c84:@CG12B?
O@-&UU-WaXL+.2=GA,@7KZ/#[gY^cdCbG@a8\QPLaLL(M+3UR&4II3)F\LeU<UCG
BN=J9HaT24([GNXNf8_5A(JHd&MNB/1SE=\U&7KVM0,3G7P22eH;@6J&N1W02,U(
M=cQ3NWXf5OL2K9B68KIc>VYa7cD(baKJEb,;_aN^RD5f<X+1UNMP;+f2+g-_J/d
6Z0]B5U086)db83<&JdM):]Bd,B;[Ka_F<+]0W>f+N0:^RWBgaaB@-FCGG=^E3N2
LW(@6N#7VC>Y(bU2+C\L]:E\6R<UF)OSB::cJH>C+aGFRcSQIX<TgR]R9\QVaX#_
_@TK@G&:#<FB[H@MQ&X]C2/c^=_FPg@8UG].+#Zb-H[14+TRg^Lc>T^BLP^aZC,I
>K8D)T^af<PQeTH2>]aR#[W>>E291bL0#a0,IEd=c+[^N5;DDRF4,PFMOO84F08d
4:gI,LGSQB7/Qdf)]UID(N<bN[cO<KDA=&R(dcCMH[3cFBV9\>25;Fb^gUD06EgN
<g_a9F+?&Y/#K)d2VH[UC,A(_=]QEbVWM9<6_b<3+4<(,)ACJ-BOdc-7)+W([?@2
2VAbH73f#ZbQ=)&]T/7GR\HIA,QI.55Ja\F4K4g^.FDDXbHXR]9L;S48.BcL0]R[
X#\deBBLdS_cAg@FPYA)SYN)#T6LPX19,ZTTYVULL0[8<S?30\EeQe_ICWSL/+3]
[g\;W,6BSZ?ARSPPFdT>2P0;-K#^?[cB<Q-],g4DBg9E[(02J^-GWUJZbVd9TebS
FF;OU&ENU#7H7A@A,E,dSC_/F6:c]Ocfe;P-W/9ZfZQ0WbFT)eB:4]5g[[65bB@b
F</7]+YN.YX+ZccO.dW#Nd7cK0ZS\\VNZ;GC]H)3dd7Q/\&I-3<YKFIY^5;M:9UF
21dYBWUNb-Vc>A1]=,XN(RcKU4bB0NAKD\e0M(<]I:1UXeA[3#1Xf@:c=R2O6Mc:
S8SK00N-J,Hd)M\Z:5KODc1V<eA8:VTf#3PN4+VZB4.U[(f-XT3UJ]U=M&M&K4,V
=^=(-,Hg?3=S>WaG^EX&H/>e53Q5S,CX4YgE_YC).LbLSP9J4>OK7=WAgJT9JXgg
^2S4bY[.EBA;OV3IE64fL6M/&Q&0IASA[O2^3]gAJ<FT_Q@0&&311RYU<16\3+6W
\Y8THaS=6E=M;+WOO/16V&F4@a_2SWdAI]CN>[;a/:7>ETI?J&,M,H[-CGOWS5OZ
/@+)bV;Q=51ACE((+#5XQ\T)g=b9K7E)0#gZgNeY.aO,[W,R;a8=+GaN1aW^JfW-
PQQUKTM2(XZ,K974J<]TH>EL9M5Z:3X^,\<g5\>QHSgZ/3H3J2O4#_3(eagN@XRf
E2WRPFQeQL=RAfXccA]<#G>c>2;c3]6(eE>Q23X1d@8+S6V(V,XBX+)J19fLAH<I
,aXER^+^=\+//P9#g[]5_CcPX<bT(73\8)@.:\EB8(g6.<MO70ZXXMC_J0J;6(?4
W7;K.>ceG(e[1R:8F5(C6JO#[KIVJNd6I?MA1XGg]H9HCAZ0b.4Hf7#bCC-_D]V;
LED28N-EK#Z?dANR6PKQ-bX23e[=EBL^[7PN7S&]DW<^21@LfW-a^:]Q?fUEXU3^
0X:)//D6TS<@M4a)^7SM)aVBAJ4K4ZK_KJf^cbH=ZFLUbg-3@,a?8U\U0@O\91Cf
P<beObEbf6#KfBC.(Z4UEZHgU1GX+.?=+8E6LDY;@5YeAOd9XVN,_B]6C^a.H)/e
ga6W).^.WM(25bCG]ZD6M(H<_&IRZ+297W)DCa[E>E+a\-[>FLY8:(b6T0V+#)#H
c(1SBb-ALfP&]X^Q_[)J.eLD2e[.f#9b;=Vb=(17,0J)9<eOa3FFB[@AK?B<CaY)
MG\>I&Q.^<J)PdT#)dR?3&A@XH,@\\+5YDV0];7(9:I_MZ/OYb&7AdBH&@db-QC]
90PH6.1S6eKL<<g?/LY]f/NGT&8eRgKf-JR#Y,HBWf0@VKEILIT&bG<>7TJ#4a&Y
f\GO@gdC@>5YZ9KR3<V#)b=G,.gMeY=VP3HOf_?Y1LP.5g?FHEDWf)Q.MIL1&gCJ
PCIK8AO@V>c)T/?FX4/_.3_dc#Jde=a5CZ^U[X,RD[2BC#<0\DeBA2Ye]KBVB/DM
-+>5V915VcIE/K^gVCa<:X7fSQTPcDXY]0_B[:PINT<)GF/(bK==YDgE^.Za^,&E
HbW[)VLY689D+LICc9FZK[d736e-XR=g10GfBGgc-E[G7=5YHN#N):S#EK>SHbX.
VTW4Y+N#5&OZ_DJ1GB<VBHZg#P(f,bPc&^A>Cd(cKXTN@\OS(H&34\bVH/F2<@^0
F4^K&W8:SM@G,N__/J/Yb\WGSb8I8]=U+=H@R8FOcg\efH[VAfC;C-.Xb]?KEGb7
Z:N_<#@V,d@WXSc;IET1eIM@+XfPTLcM9U,;I3I9+c/eS-Z<Xe/PB]-#N/4/e80;
LPVON#0:S-eE,(BG>/ZKc?AFMK,G4^:af[Ld1Z7_7_SS\)4<^],KbDGK/K..BD?B
=&^)06\ePfMWV1@F-0=2/]1TO5_AeDf2CKJKSRAg&;CeZVeG]acUMTMAV4Sbg4JG
K.2DB5-GaX&C7Y_3Z35?36VC.?ZbTVR9_dK1#VfXc.B&95)?M=3HV?#.CD\6O<?L
S-?UO+e0e7PITYaE9aXE;K&MLbG@R_Oeg)+9#@;IH7<\Z:30)4DM#SGGY2:25-cb
&C^95[KZ,@WW/(#3J3(g6>5g)2V)/&8K0d1G#Gd;cA384,8ZMJ>/J0H8YA/1Q+J^
GfD4HOQ>BCFBgb,2dCFQ1:T+27S6N68YS/4bcIS(?FX?R3)a-e&d55A<94^CZ1PU
XTU2eSCGFK5O>S7J;X^9)+D0Pea[eO-PX8eTOXEa,@^4;ZM[bGADQ?POIM\]Sb&C
39\_+E-H0b=8#79OZAY]8M^535Y3;]3&B:RJ>MN:cLXa_FV+c._7ROGF.THL)a]V
C/ccGDQ6K)OL^VY[8?4Sb>P5:T(R-IIX_1[aCRN4>;7;K&^7EZHUTI]6DNUTW0YQ
<M_23HZ(J]1U9-AP)B-WgP(^T#DT^&d+_fM?(C8\+Ta5QcE=A>-5f4^6<-+,3V@G
?bM?N26(Y.U[[S,K@T^VD__#/5)3^gR<9=/J[^9A[H>R?)>&0cMg)82\SM8^EUa<
_B7A#?0(5\?4<a5c&B3bd08AU-f2S=a,MTU+#6Aa\5TMgLE5^=@TJ)Y^=TC)Zd0d
:TLO,;/V^H;D49X]CbAcF^#HOTC3<&#(+,<eJBW=5=\f329_5V2GMd>-+J)[BdFD
],3ETF5+=M)6NR)>AQgc)_dQO:(LP<Y82a)9:FSJ\Lb8f;&^V@2\M]E:d_@;2A??
,4Df+1_))7a=2#SK5O>V.dL;Ia&]\F8MR?f/>a7fKaDG=\/EN^[=_0_[[9-4eIS@
\^YTQO4_G;WNXDTE[:\5[FNCZe;EJ-Lc[F]@<ZefQJE3>?^5,7/_-F+B:ECUK[f4
38>:)V&AK7(/4[9MUJHBb6Y1=PSaR2(Ud?&Y2M;C?PHLeMK17/32Q^U#ZA7XDMeg
cZ@>CJUW:=\H\BaMY.2d=2aGP/3BZLOM)+)d:FHG&.M6(M6P3]4H@MO^57A2S1^4
2,9(L18#Xf6a#cEbc;I^PAc]<1)/.7?JG]ZK.d<dP37ROCP\4e=c;2a&bO[55TXa
H>@U^5KZ2^9/M#2VN.a43]a7<QZbP;Ca4d@]8Y)\=L2WH6S>=2M;N+CX]I&@72?4
1QabXcce:E9XBY\,U0T7K]U7S38/dR?<@\gd+N6->@AYVH3TO9>Ye/8/91F2P->>
><c_<9,AH?Q9&b5X;>G^^H#WDP)8,O50ME(RA=\M=TKH[6?T^(1?@H8dP_ZT1\aI
5,+98E(LKZ+X?SXY34La/TRT5\RT]2a-Uc1ACK:XDe?:F]XT5-1EfF([[A8-CFT2
QMYRG].GLD#-L6)[F_T4PeI].,5+:B.E_,1TQKe99:8cJ\;FW-LOHe8)5-;PW8?2
^ZR#7^,Fg.<_=cG-/_[B/[+U5-X::)#37[UT,Ie2G7:4L>1GD&N;5cY^;;e(.2UH
LR^0^AH\OaAS<+_[fU:9,SNS?,WeE7Yb+]FDfUecc2TRB_V3+#)bSGW,[<?Z^TWN
7&C?JCC-(G8&Qc2Z<cA1NCK[SW5JAdAQDWS<=W,6SI-/Bf?PaDHSH0L;)MD9.Hg<
)#_-;UYf(DDP,HJe()7L;JCUZME^L;>;PA7KH5BI_R<0)+3>G6VPcAWH@QU^VDZL
\K6@NN5CY:461KZSZI:K?KQ.Z^#Y>?73Ec&cbC1If\-:gP6f2Ce2KW7^7;SN6GSb
&HeBNB\<\S9?JZ((>84+[PZ)RIY6[6U==gQAUL/SS9bEGARg^e\4XFO.C#&730TB
G=U3)SZ8K_gG\-KS2T0--<+J[SP1[JBJRSKNUd+>5YUWc]&G15R0>(^<g0Za.HC.
-a:JgX\MAfX9&5TONE+-5,+I.8K[X>AZSLA?WeZU3UY.aKDaWa00&SH?\(GJG^P/
O,g3XD8-.faAF<1;PO.aXY#AFKWDe?g[50-V&d\?V=BQFd3C2WC6UOTT4:Sc=B3]
[1ZDaP2^NKF>2T0P,K1-Oe;)2V5LREgN:Z+I[H\OOLb9U4J3PAI>YdeB,2<4-90_
.Da0<abNab5Q<?aZ.T7W63+(H+R)HRbebZ<E>18(YNf@UC/a>Vae90cM(F6Yb^:I
Z/6Z47gSXI(2@+I2FA&B[N5d1DQFeU6P\=Yd_Z.+R.<XEE65_IHQQYLf-8cA6P[3
=OENQ,.E-1\PU&P]fXX#..9D+4>\[,PJ<ZVGLPDD/CgPG>MeG-;;\8QOW)WS.ab]
E5QKS+Sf<=NFg.PAH:#dXE5ab9)_8AO_E,>SS27M;GISdFa>CVGb.T1?@0FBL.BD
f/G_H@W[U5&NNU-2OeAZS/UQJ12X/L#@>5N9[(H/,F5\M&QbU<U^>gL\\EHEfW73
QE[R#1g+W[3;Q1&b1QM[\La_35@bV=<gSEJGK;,bSLcG>[XYe<eLGb/R3Zd.C6QO
;;RL4^B=3gaW..;CD5+,Zd-E(;-^:\>?X<Q[MAFU\&@5V?_<;DI#H30UT9^J+9fP
d,W^6S5M7]03<U(/YWaZ9[KBZMIRcb5U\HcERVcJ]=?3_BE#717^18W@=C^H^IEN
G][/NX^HGE[C+-0_=NFIcaRES1/JX?K;aY3LJ^+>eWCE]Nd:NMB,XR=34(0N@&P:
XFCL[4:G5O/IS5K:,3d)K?8B(cO,(R?)6_?HafED7M@ZKYEB]TS?2(CUD+@N_2^P
V1DCJQVEFQ52UL6bTF8X0(_.6Qad&-KGT192-SF5DBJ/F.\755C/Xf9#^KT1a3Y]
-49FAOg@=&Sc+dd?_E@_g=8Q&?J(Ja6T5TbE2@@B?[AN.7EF,gA+CF(3DEg4M4Q:
+8@Pc(\;<YNIA.aYe,:a8U.dPP(#0):/&]Jb2M(EH/1OJc\gWfMN5Q0VA6DXZd4[
c;T&6A8F<A/2G8O4f<c,W[P3I#_PQ@4:K6FT&:^AbS--@b;UfYMBU?NR]<de1(02
QU@.aSP-Q&?/b+YfGeg_6CSNR&02a[]B-S>JD[bLV/-)&=e_;=aNT_]_\dag7,;C
Y_.YN>F^N/Jb=_RCZTYQ#JTBS^WIdP\Jge>\),K]LTaY&(MMBZ2E<=_PVWZ@>,;A
MXF6.[Rf/D7d7GO&32P@VZ]?\E?.ZZ=6(<+P+Z<&0<+P^7WT2b8DD2;@&e9=gT.J
/?[fI5>\+FR(?Y#0a[GSeLUW,U5C4gC?]4E>07eA@_cE85K1J6f\Y]ObPb+,0_-_
5/T1(;UI1-DD4gW[8b,Za,H:MTWAM([e>1e(g1=\Vb)aZX)7fa0,>bIe@7a&YRAQ
157].^daC.^?YRG[d8W9fK3+5CQ-a_].A+2K:[B5:cV<_#.@CGP>+ZH[XUB7(1e>
YV6?c8M^O59@37L^2HWFLQXMAX1#d;)GILW56a0;V94>cS248+SX;LPU4:.H>;/I
O;F=&GSKIB&De(.96fdG1RRK\&>?X/OKV>,(-0PB:Q6544>R_KE)Y-YAVX,MCVW6
1fMBeg?a?>W;e6M.d:L_:Cb@11[^f2GLIg7f9Vd0N/Kg7+7Z)ZXg4\B[GXeeZ&5J
JD7<Q2J/7/eM7<:?eWI@ST5^gcX1a55[-P#X-343fE0.#R.=#,,Z#cJ.)dONYe1E
fdXaM3I5^4;62(_[@X8JH+g?1T:;c^HV.Zb<bXCI<cbgEX:KT9M;L,fgGU^JTI(]
[cCP?P)G[g+6BP:G>6e6RA38<>@fMQ:/CT-2=2fGHU._2EEWYP#-0:1\>-M]8XAS
^#K1CRNIY#M1?=7RJe[2;_(WfCd[[)W1Z(V:@=4RA2g?IfWZaSG>g:AP)^YHD:cE
S-Y7+dd#J=E/ZUWdQ/N:2S;HFPgVX-CY=;(CU+B8]BF;,Ka2+5V)4,\+<-S^S+\S
N.=6)eZ-.64G7(_8/J?H00;d/4H+c;<aDK\6Y56.N5c<]/;DIH:fbO)>bYUVK&4P
g3W)gZVgROYd/#1R->AJ3?A&6O>Z=@);OfI\-7,]-H:M:Yc^b2U.PQPMZ9_\9U#(
RNKTB0AUecJ9<Gc/BI]KD+cT=5]g?ERa<0R1K[&NaS,B+YVJ[3DNG:Yg\??YfHDP
=I\CBVCAZfQPa:d/e7Q436)TG]77-WBB(MDG8dNOA@@9+9a=8cVD5ONPB?V3?R:^
.@N,D3Y\//K,-OLS&)0OJL<_ZH+MQ_NHM_E,Xd-f2L]PO;JSRD(5@[+2-X-+,e/J
WC_4cY-DbY0:IAO\2607@:\&=dC@XG5bHKYfI8)_T9NaHN82f_.L]HfNf<]:Y0Ec
1K:9EM[24KIOXLOg<U;c0CZ?<+&VLa\K#U73CS3E9aS0a,<ZS;EMQY\]a9X4SZL/
5Z>R5C:Q(I_^H7cfO0RJH(7YfCNRO#]OJZX#[->7O3W#8)^AMFA0I09X>Z+5.V#C
fMV&77W7KM8#=ce0P:,Lb:ecI:G+>3]AQ)UDVO7:;&_YTH>9c&+fG:TO==#geE9K
R8HAN[Ded:>J:,C1BXTa7U1C.M#N#8#C84)eOLTf)M8_AL?4)#?ScbS(KY0gNXL_
C4J5TN>[GP6.T1Q99;P=9d0X;N#(-5=4;HgC/W;@7)Q3JH=^I&X./GY=-cNUR#M0
<8]4:&VCP4&\fJ#aY@V9?eTKR75/0ceA6=D-_5V^3+.^#B@HJLYFR,K2X[563=1-
3<=d1=/=\a:FW-2IVA+##YICb\KagF\Hg&97(_[:@3G6O\MTG&2#=6+L)e?Q.4W1
3g[N;C@8\A6#+/3d,XdAT#YIFKOF_ZA7cP?0gOSFe=9@Ve4dBaJHU/d]Be.<Z]a_
..QK_09W\TTVUWTK0..#)ZNf3gbaA.^JQaW=Ud30g4aR&S1Q##F8F)WW4:Q,L]GV
5;abc/6^4B929fF06C9+a_f)U9XX8=P]E8#@XT7[/R8AZQ4?DWIYD6OG\GK)#_-2
a8L&@OQR/DP8ZODWU1@H41eR\(KOX>\F9cg8YQ^A5ZKTP;CDLJ80C49M)]W]:5QN
,R[DGIRVI8Cd>-:1.ET>37dUJa,FO7A1SbPE.^56HdZdY[@T(=>GC@36@U/1V;MM
d-3cb6-g100V4BF8]#+=R2>Rbg@]J_&N0:b4g97)\SDO0g9NOYI;S8_DM]O([?4[
NUU\MW.U\D0E@4A+&6++gY.DR+AV3O5J\E-0dDD4@X=OC(A)^dDQ>]W\eTTPfKg)
Hf&T>7C;(/]K2X]dEb,Qe-@36P1U>.gPcUKEOV,H:e@8++^AVNJE/]?PDVd]==c0
JFbGUdJ>]7E:()c/J6Ld=F^EWH\,U&da4:eCR99U@SYOFWW9D#&=NZ5TNL-ICXc6
QKbPaT?BcONgI:9]Ne\;>J12AD^M[bE9E4/L&Hf?Ec@G,6AgPE5_Q1=(9DdWaNA?
cGe=1d\S#Z5YTR/f6S.\JdYc]UR&eRPfe:fHD,J4:^1VRTGKFD_G[MX^f9R3&+ea
e8_V_#=eMY5/DNg#^#)JR8ab)W6+1^c18dD-?dDa^K[5_b=WAUe_fKb8HJ#:2Y^>
TZC=)@GeHQ8BO<I(YX&5_U5H3KA]_1DNb__]EG_b,Ea(e[Y9]MWQU1-FFL_<ab;g
5VF^bH484XC)&Y1R\aNQ;L;)9;@,@b(4Y8cV)=@_\K,D&CYTg,<R5RYX/L-b:9P;
5>TJMI2@ANM3-^U7?C4U#.;D_d;S>[T/:1A74KcdX9\M5)bL;U39MaJ<0ZZ_0XQf
PMYPSWV@Y@78AV/0.2IfRQbH96C6D+JYNTCHV@35F\U?MB.6aC<B=a,P81Q((N>M
cCF_E9Le?0(\D_M6\^Fa4;?Me;CeB._?ERD._N0IFUBe@I;:=__Q>2EdBN(+OWId
K_54DLc@-;6-,6aOESO4f<,??Va?Q(;;;1R>[N<[4]];D)CZ#+;V#b3.>(fM<GZ_
bgP9Z^28O&HK#9+A.E[=MN_ZBO\)aDNcTEE;e_GY-ScJ#DF.-gD7J+/4g6X#97<N
RNLQ7MLH&BP#B\e8_fIX>8T5KX.Z]+@O1&XH__f)&P(-(9+>9AH.82+R><PGAaJW
1>0]^>E?L0+:e_Ef^.?=f\LAEg6MO<f^C9OCR2bAVX(PSTS=fUZ>ZT[P>=1+24]6
Z)_7d7RQb\XaA=aFa)DaVQ1/Y0d<:,DX719;ON^;g^6V8;H?@;=c\]F1P2HB1K83
=U7YWGRY3(V_eU;Z(M7VP<FLVNbJQ4F3?V)-Deff(8ORQQ;=Z/^<7[Q:T/c(gF8Q
VLVWNNO<>VEcC(?6Xg(e:>\MDC+Qc?NEZX=>WU:.9OgHC5YE8J\T:CRe):[_,72b
I67UTbbNA[T=)6AG1bQ=\ZeBI^[#4GWC,M/<d+8?AKI>TMa1#A6VBb>T7Qd==SZ-
-XAaJ3F:[DPYBUH3//NLaG#abN^J/fZ+cK:Q,LcF\f@#OFR1K&[:YFB.C5B.;8#I
g6\OXVc+;96;#13e@XH7Z5TRa1:1M=b\55T+.bLKf/e?HaS6)2GMcJM4#@Yf93FI
47S@>=a>I+(O91?c7P3\0dF[4\21[FXOPE=\)>-,?BB>ODK2#]EM,GI[S7\G,g20
8]^BC>D>DP(LE12BfGgg)J,b<-4,-TB&@05K>_-Kf:)9JP.O7XL,6<C[KceK6CBB
J;8E]>)^D4U+=Z1L;E;1W/08?25L,W2]g<IS]ZcJbU<#6B1QV,XFa#\@>BbMD?R1
?G6CdN7^Ng)+7/:3@>d\T4)b8Sd5d;2HfP7M-T0G7[c_ddLL(8)>^Mag(;G\EB+=
:WHJJDX&LgX;/b&^R\WEL(7TTg#\;+3@--]>XXg3EY=)B=YEO=4.DU[XJE3T,RXK
Y<a-Q-a(=YYc?[&JP./&bFQf)>16MCS[W95<ZLHH62978AI:C7CB3&SX?1#gSIT?
Zb[FCR@WX4R>EQ:=A09]5eU8KU=R??Yf?&0Z3[fWH^<J>B8F;L\d=a5B)^e<b51E
RcLVNNGDFT@(XHO0b+/R2WO&,R9U)=G6V_f9I)WS.\X1fM3.GX95_1OMKW8_F3AH
U<UCUILBKSU.M98/0)(AZ9)72;FEd:U;-\J.dEXQQP+AEY_KZ8<<CS^AA:>#=/T,
D??L#@f4_ZA3aVA8T<b(>RWCBaN6Q=0TX#\+GAQM9]9cXJ@Z9OO6,CJ]FFaTHd87
+ZNd2ZA:U3FeYOR-aM][9.5Z;;A]0/Y3/Hf:7V-Nd;0@\^MHcgSO2PE=a]7=E4D7
g4&cG><fQc(BW8IVSY&HH=:a9gEJNIUgS/5=WX.MYFa+T;PJ:S^\Y]FT1I1Vd3FZ
\G;.)5f=Q.+1G\/>?72]c3LdcN9/]\[^^Y(ZT((01XTVR2)M=Ud4L@[Y74XI<&IT
cfA<YUaPea^f0@(#RIA>.B-[>])0@:&8Y,,GDB2)9GZ9a&>ZBX<+UQ=G2P&;V+BN
?@V2C^(P828dbBS#^UPcI0N][-I3#=3&6D2/)FAc)JKT&^G;?2+TT?D8#_)_OXQ_
Z;]b]-aGT#.gGeXJ_IZU&LJMe=BWdN0O=&F+.a#G-_#:J7W,E-IJ[;VML5/cC,B8
YAQAHPeH4L_0FJH.<7ND\R(I_KT:T01[7ge#b(2-:Y6\F--HSZcFET^N2/P&3cg,
[:]I)X2-Z1X8;Y#-geXDM=A<YWEIQ,61H7X3>-XKZS7UQ=;#R=dg_:Y,?UL2PW36
be;3d?dS9U.[cZ&gDBFK?^<2dKWZ\-E8A&;62((bQ:;&Id/G)F+_ac9>YOLY\Z,[
&:,8GfTeT8[4C](a>6=-VYBa3[S33K\HEdH;b==2990K7U(GAI>9aDe4HM^6EJLY
N\@/4-:CE5;7@4I(D4/\bd-dJ<@(\G64YPR:M09<=U/gfWE,>Hb:&<YW>4#IeGS#
73Lbb(R/].d&?dGVAe2T(>eS663AB7,QKY]QbC1-#cIRK5/CG1H;H4=<4O=GFI^9
D#(M67@=L<EX[RWW1fY2OKdI6=,cSdHEeF9W[,OfK>]Z>R0eC0TP1a/CYQ9PeOg\
e@GE2Td1[N8E3D=83,WEFf@3YFC.f=D)Bfa38Mc+c#?a?8P]T.(P>RSZd2Fb(.M0
70<^WW^GZAXNb-WG-(/#_R3Nf]XSPGaP<.)8/?I64\-OQ\cK>)D)D_]@(?UL<Ubc
d1IA0H81Gd.\Q:7YV\B7+H/Q^QQL^.VGMIT<gF?_)RGY4NP1OBD6B2Z>;<Me[:RI
8(O9F[C5U87N&MM\<;\N,UA&.ABV:ATI0,;QP(egZT4V-O8++7fHCEICOY:4S\E\
+#fS,/7+)B1@?SEXZ,E#(MRYQ&LD^gD8B0&cF>5gZ81d,Cd<AQ9=f\TE>@9C<1fF
bZEc3?B7OT#Y/>#2C7Z<JCf:]R8:GD@PBSB5-e:<KARZ(;L-.]8N/g(8YAQ\A5=?
Zda27].@7C<#KF5/^#R(5.S24HQYWaS<&DOH,.])H:Y;BD[V?;OWFM8CadLW]>B/
)35<328BBW]RFQX@M+R5NNFPSBT84-^79195_J>RbR)Z5TC6@\3@;XM3#K\</a;_
fJA?_8Ld<];cg0^0<>0[C=9X-Sbd;8MVa5gBJ0)F5g>978ebT0^I\G?6M#DT]WD[
gI/e](O@DZCM55V#]6:20)J^TgT7;S5caX>2_6/W\033HHK(5E]D_+F.#;9R5ceb
f[T&=.D-MWQ6D+Rc51]5NYf+RcaA6X)a6(HGGEJ0=.B\29([&G3>X3KUT>9&E[Aa
S>;cY3P0Af@5M1881a4AbP+1D#)I]Oe2WdB3+-P37R3V;-L@8a#-B0Q<+fUUS/cG
HU@:IL@SGC\0O_7U\-#KOa+NMS\+;3#Y&.5,5/_ECTP_Cb7CW(>#?R[NGBd.THX,
S[aWP?JPY/4RgX.#7H;R5S3]V(EV.RcCG0.d+9?L<4.98.8<a9E4OFF243G>I:48
N63;.Y0]FR900FHfYQRda7AH;09EGgQ6aZ>Y@R,<c>+Z9]C+T]T7d]aEW0^#>R79
-.S&VI8E4VJMGTXbR#/1LHg(;.H,5_3JWeB)&-GUQ&N[Xc\U_LD@9FWFZ#/CfN9-
:##6_0GTR9F^^[d^>M<<1T)Ub4[.aN/Ed6dE;L#5XYOY)80[P?F]aJ_AJW0g>;E1
NQSQT#:9XNB9NG)39N7I8,X]2[JNLEeaELQDRc4:.>6KYD(B/GSPKD,^<N3GTOd9
)S@)R&UCWAHQ)T<675b-:BL]JJG=(>]cUK<JgBWJJXMXGDIUA)2S;;[MQ322TL_0
.+5)+:)Vgb<<5N]^;+f&@e<OVg0RTR>;M);,2I>^&,5]G8A=D3AH0PC:A)OdS911
RgX_YLDU2cO5<&H2Z<COMV=M,7XU]fC0IVW0LJ7FM/WLL4GdcebLe(QHI#2?[e2Y
.CcSg6#]FV6SBP3aC^V,DAW3A;Db6>S\:?)XR3]5,6a;5CRHK04XadSKR=DXEU&e
F/^;;WQA>]#eB^,b]2&H<4]HE>S,K/\9Z9H&@AXWK(.E)26UN(G9&3(S1^X&6#dF
+,4,gc4a0D.dQdI6WaCTd2X0LGBb09+ZOBUf5HNYL1ES>ME<JEW1^F@=0(bX57#M
FP-J0P;E1095CaX]GO2E=Y1>KJTX;EbDKH@a)@M:T#++&HCI[9YCKHC#<8aFUgfc
&0(H@S.&aA5[/O-f.T;Yb:@a1e(XZG\14>Y>G<6F&-XFS)EY-aALD<=R[VX8G=+F
ML87;G3a=-<gG.V2.dL98F4JHN)52IC9VNR._&D<B@573fB>db?^._]R^>[J,8U]
9?\f01=[f;R/>:\5>K4Hd2]_RD,_-1@R0^S;cUP?0\SMCACZOJc=KZ<a,ae=+]KD
Q,c^.T>1U,:.e]9NYD_0_Ld@?>3bf;M1eR6g;^8A)JUF,?KHcQL.3HIZFQQ2=#.K
MM]WRE3(Tc2Ze/ZP-]]1GY6#C0cgK1d5^?<(=]4Q&,R(MI8D4VPJC[eQ7Q.cLQSN
67Z2O&RQR]d6#?36SCb8G6DWN6B;1K:OV2CU8F.L:W@>5@R++L[g.\C]OHVIMU31
VQ<MDV5#)edG+6+&B+L/^H9:F:E]O@^(6=KRY24?cU8RN3I<O7d5I7KJ^&NHNT>;
:5?7eW9Tea+[QCaad2cBAIPd;G>CTCd4^ZEJ=97:C/].fg,F:;C,D#a(=L74^I>6
:G03L7N^?3;]&G\VBB\RO;@&B;03Z=?5JC2G=_+&.7,:IJR(&F8NcVU)]:1R7S+c
dD#7;_dO5PE^CHPWBQHC7Oe:-W^6[Y2]Ab7B)Te^2QZDg9d.O,2M#^HA;&BZL&_I
3D6/ATM@1[::4+BGT_.:YBa>G<B8cM[X5P.Kde\I=eaJE=ZZHB750FD.BF9ZEZ29
7Sc.+7H2]>8/TF=E=TV?R9JN1T8]0KF\c[U^;6;18P4?/1-]C1f?=\XdIaV2Vc)9
JJ:0E\WSS#]D.)a]UMC7S(V0+d->&GUJJ=R_M97-=73+C44>6T.AQ\/#Y65.f2/H
V7TIU)6AYY/UabEQEWYMM#02]/A/<T1K>Z4J;34a(66);/dbZf&&[7A/+[-IOLDT
+2/P2N7A0G?0X]F8R^]Y@MNgf87UaO&\EI1[HC[:V\=g&(+TMW7M]B<Mg/3,ATg_
@T\TfIb=F<E-?a8[.73-A<U\A6+1,5I5Q?R=(5PKT&3#+8-P5N]3X]EUc&HXX)Hg
+8WZ</\MBXB>92Y]D+BbEOUB6]<T0\4gA>Ge&G-6c.=c@OS\O\O+U#1AN#VCD[46
HcKLL4<9_bSWE+Aa^Y6JI[/Q+dI9XC0J[CZZ2D19_[Da,+[Ef^91aKGI6g=B?.36
F8:bMF3LL<]Y)F:@S7+DUYL\>1M-0[)7gQT[NP4/P]04XL?eeY^RD=9[]b)@R8Y2
<:P/2PaO?RE#Y7&<2<5&>J/fC8I3ER)20T5D3GFR=6KQ2^e@DN1BYfZOY#_7[_5P
f&->9K5Ge3Rc(2eCGZ0I:_gNIf3;abd7DZ5J7<#(N<6H#(&+QJ=.6+E2[A57D710
=BJ2Z8@;U_Rf#ff0_O8/eV:B<([@0AEYQdB5,^UcN16(E/]c6SV49--Gbd>6?MB>
?KLYNa1_e+ME#FFeS+b_e(M4H--f^[MEFR9gUGHM,UM=Y#V4a).TF+Z^60R.=MCd
g2&]/;,\,+(aR^QPRI11,_]SYDMF3X8XP?gG.1&BZDO6eVb.ac^)8C4a(R6UFC@H
g#7/\#.;IT@=3?6Eb2F&Tb#<HZ.]I0&?MMT]9.=.FQFe\5@M@H1L4();BI[?S@)a
IG^ZbBDa4ZDVd03=V=.bI<LfD3]^=O0ga7HR[M6QM;(-<8<fdA]U5NJ9=@S=J+0c
:J6T88c_]=Gb2G>FICC/]8QG#+cVIfB2&Fa[>0&(:1:>ge2bUQFa+UQ?/e0(.MW@
cPDZ^J)]g=W=JDMea-7FYP[/gY9UeOe2.8ERQ)GR;:;J:]#f;BO-a(P48#3^TYF6
6RL+Y1]-Vc;LO2[H?C,(MT#IVS::?Fd8QR)CJGA62D+7ZDBR)a(.04]bPaXe/)D8
,4^@4&BOL@(SF9,V;-.&Lf5]?3(3E-(M]S(T2,_Zd+:A9gfCX:X55gDZFLNU;d@P
c#YN3VV<Nf=d+_/3<;@<c/d[Q0We5Pc-33O[Nd]@KYg\DA9+,7@ZKc+5fMOFWPJK
_9EN)aU692@bL#V24:W6,.KUc#&V]Z.O-CQE&FCI@6YC2b);EbH>=?E>ed/fG9@:
:e/Y,HeRcTSbP>>N5b@Q:+X4P&OB@W=9ZP.==/@][.U?3(eeI<\LJ)C5,L[IGH6S
LY:;&TE:3(f4XE1=9g7XGIGa-6@1JUYBQHf2.POOC4><GS,]5XY@(6RFW;Z=1g6J
3OENe];>E8KI0)[?L2>WCQOC/Q&0R25c@E]QGeIg..[fL?AfLe44FeWYA84^MMM(
2NbI0)c<58C?3T^]eC,+^&@.WG;L/S=@57BEBUN=bF]Mg;P\;ML+MPF7?/5N#.&+
abV\9fC5.IJfd1<JOb9:AYBGKSVbA(WgVaBdS4AFLD@KPQ<]ANP26&?=YLP6Q,dM
/ZDFD7=87)+^0[(#234@;BBD@3T->2O[<^[+S.-6K8=YfL\P:1[:45(c(<BOY97b
bbc.9#dP<SY4J]8d:)EY:g;>J<PaFHSREU/f.XJ)-E+.aMdGSR]:[N6L2>^Xc-9B
3/)-f@C?dg+>SRY/1Q6?@?X\Q1N:ZK_]/Y1KCEa2cMdP/LQV&5Y]gMUAaXde9;ZJ
\0/&<NO>A_SAB1-VB<b+^\R2V>I3gBZMVUc(bHIP@e)E<bU>-)AaB\L26dL4#82]
U2433D;O13_#ZA=7c6#^3Ib-X.XGS?c=QPA?gdZc>35#(Q:HEAQ##IHLY>,eYefg
@<96a)8PNODI[PG(;9e:HT[.6_MN]UAfL-H>a]X8YK/-84TY)OGagFH8R_8.\2Ug
J)@N;N#K>7AEbJ?]1]@H]^EfFNS)\NBEI^8LaO>?A#,YFPT,e52:b@=58)>)[5Tb
QDL>#HMGEZ6F/C1(C:Ja-\.TX6A7??B^9cd;^.)XD05?;JCJ]UQ?gC6VSZC.5:[b
<d<7W==>,3DL7&KgI]f6a+(8B,[&]Z;>I,]FPMK]52W1J1_^fN7ZSM0EQW26#cfL
MQ/HD6a\@f.54YPVP98E:.DOU=2db/0^YJB8.X-,WJ0^^T(4a849@(gaDPUc(^9H
ERP5^(JS4](6;H@6?]-Y:?fg558IY3^bVM<NM3/2Va9)^ggcFM;<:WHR;KFJLJ5[
e48D7[CYC1QefPOKNN/6bKJ>ef@7J-G;5WY6IR]CBV,8VR:J7\#[2.EgDcYLK1,M
BHFVe6QM?HYDd55@01@.1R@WfP4B3=3D-Tb8Y1(7)3c24_eI[R8_;cFN(H@-db>e
S7Hd?AL6L)XHW(:.&_J]3LDY+QPcf<IcT2+e[:AcKdR4K/c1TT1[]J69L)S&2QFB
\/MPVFF6Se#dPg@)SZf;[7@e2-/4W)K^?N[a/G,()6FG:;-&ON>fT<[Zd<;)Qe6P
WUA[EfKAV9(<Z2^[&6QW;C.ReUVdT-NWc.1S_#CP5QZV;775<Z[91C5UFML->a2-
=E1?3D-E->);aTYX\G(U^TFcI4gM8P8b@;Ig2\T>)T@^bYb+d[ZV</X:a1RT3CSY
<\,:77JQ^;&<702(PPIIFAK5^UJY5]&38?,AegAa-aLF9[aOHORc,(>RbaPC1g\+
;0P?E)&)e;20LCUL^1GgZ[J4176+/X)4I-^;d0-(]<>KORU&b,]WX=2(e?AT6Q5,
cfN\\(PF4cW=3XYNb1UF=(b>74FUgf6gX109<O<T92GO>H@U@fS7eLg[?&<_VQ<J
UNHT\T-P^TL)^K@?cA8FLDg_Q_R/(7RZ+&6QMHHM.J,9V/Xb?G\:?C78H/42AgTI
0=OK8D/WVBXfG5>DA.U\(W1TYJ4O<(@f-)U8bQ(O=X;:fF?Gg?B-dV@NN]L/1d]+
L0K&d&EPN#A2\R\[PYcGGH;@^OT1/^&=fUc+.74(IZ8;SX7:N&;3QJ;X/Xe-X-gN
NFT4A,^QKaX0G01MU9Z\)5DefETL\[FNF5],aEQYfe<M41<^BOAg&6L=WHV\<D5V
CCSZ?CT2GT02STKA<0d+e(X\R4@2+O3]Y\MX<gY^f.>_UQ=Y;]@<0A^@(D0UF65L
X-g)d7VaM;ea?PK/7V46R=71c?3JX\CLT;-E)&Y7N?Bc45)/gG@=_?1gT]QM?[9=
Q-67_gEddJW8WO]1Y?K)g_7DJdI.4YVg9ZM4dVb)L:e#LXO[5D&I\/&=Q8a@.9Md
[LS9);A/<RMN]b=YN-1D8BK&],^.0?RG\_(N2B+6g8.C39^N_1-O1&JdJ7RGYLe4
@4(ZEf2#cUZ(_FdJ9:[J)ZYXMa+[<K&RO:=H=-X<Z1CLf4F9:VF7Y>&=65_=#UA>
LW\Cb2^?^F-3/:TD1P_LA_;FU>6_a0D\(M;:MZB5IFBMab]?:96A_R4V?2a)/BWD
,>RB[#22DU912\O(J:DVg;]]Q0WW[@Y\:;a.DYQBV,-CG>000VfS2UgdC>?3ZW6L
LF(A2E-W1&3,&[b5\IR>]R..LOU]P9]3bRTRT4b/Uf955BCG/[05?>2KI6HQ,gb<
C?fIV5_[ge-_QfJ[2P[HgXA>8Q/#gG0Sa#=,:_eLgb8VR_b<]bLW1XVJW;SOC-_5
/9b5TKU][YL+DgC=KZMBWWA,C^)4^J^d#XA8WQNg6F83f>N?@):C?Z3dY34;<^7g
bF:3d90NgCC47g0UegC8,BIE)=0X;J>3ac1g:C9:WJBK1cO.Xc0^d9GO,.30cOXB
XJ.Q7I@#=;#<48T0S^]#aR4)1L&Y2IKW7,)LTJG\9c,GE5BFg8JL_FXb:2f:G>6R
1^=-8f7&7X7_.GO82d))(3\FK=DEMY4+&5N<90=:H7_+_]4)^+VS92QV+YPKcH_]
J:DT9-=?2QU(@BO2g2#18_/aKZR5g1-1HT(g-)-=HZ^BUK0_8,@BW4?JBB2gUL=+
KO^.=)W1GA(?\XdNgB?+59&FJQNcG8)8;9X>Z#4AKcFd4#:.-ZCPM5Jc)IMB\;R,
>@0f^R&O-YH&2gD<Pf5ACUCPe;A6)KM2G<OGAA6POGMME\WG-)JCK0Fd<_70_6M]
QH9&4\0c84E7N&L_Q951BY[UDV.=RgedE0&g1=@V;XC^];FJR9UL\)1&3031YaA?
N7?UgQ[FIG-VWEg>fGM+85CL^f]?/Y2[NfZgAJbEg301U&5(&FO@6D;Q0??->19b
5\,a@@V;M:#,cUSP[28/KDfFGBfd85H7eCVUd6M.FIBM_HP2OS6:>[dFJgbUI.+f
@D7C<R0:M/W=7>5.T[B:NF^RMWGSXU8gZOG+?b8KD.4)BD3d1<1cfC3R5:==P3DU
KTTQ>H8KX\,]KK<BbY6/b2eNVcG+(2Ia0&XQEH5U/HXHGee^BWT)L:CRB#T;eXW,
;U&6X33S@0:HAI;FP#3d1KP7;^L_e[:LCMgLHF]T#=cK:cf:feddW_B?D.58\1&T
\R(/K^.L=PFbN=)\(J#I3.d12O4Nc^](W&?4DR\W=A>>+#DQMO-<8gVeS1AD1dB)
cH9)gX[[UOAJ?9_bZZAV?TBKWPO=/8Y<5[60UZ_U:#GR#_[.L8_XDU<#8c5PBJBa
H5a<T0b]0G-<=_9=&\;(0D?+g\=7bQ9bB?STI^YaJ556D;8IO0<,Y]<.7ET)c?b+
X1HR8E5Z&=1?Z@GT^4-#9C7JKO\3]D.CD,<+?>-)8/a&BZ/SC<gF[9a3[3XR-YU0
EYWF49N==ZV/ZJERCO#Jf8f\S41=2EZP,<>V-?.\]a3gFK)&g,RL6^S1YLA0g,SQ
3C:40I8YJL0?ad&gdc^-7FQV/C&1(2]Q9QF2]XYHf5PaL:N[Ne--(FP.EZAHL_LF
O.)G#\&K/4\O)f)f^Be]WH&:Vb?Gc9S.7<H[DW@.^?,/Kcd&KC,(BJ[+&RSBg:TZ
0Q=fN,9HNPX.OA>gPg;H^@@YD#_1F#Td)9_X2U9ScfHXaRW=\;S+87X32IFWIPaO
-7-6PYE;PAfD=Q[ZZHEFVb(b^=\S+Ef)QK043[e0UU_PZH@K[WFAFP:Kf6EcG9TU
bW_0HTfQ,D@_PeA?5C)>XdD8V-A^D6?A7Y#)@SZR0H\._/FUA7=,H+74fHC8Qe8F
N23F0QC]aA>LMDPaH30.ScEI-NF.R<C2/X:Y4ME?4BNVFF9;d:=2.Q?RKHR(=f/]
d2[GR3#geaN</#F&:Q<A9>)PKTM8<?+e&)-=8WVFf?WWFAQ<f5Y;EI@(X>4^,4@S
BGQG?@[4QJ1NM5R#_.<YbF6L8@SH7[)5?23a0-)Y]04a=NI(ea/)eY-@=a_AQP(C
a7PdL2cW5Gf9Y&[YbRU]8/(W-5<43GY^DFdWGX\;PDIDX\)&CX-4I+OR@&Yb-@>@
C>d5]/80LaK]?TSb2&PaPF,P+S4g+7P8RH#HEJ\A6<..N\N<aRf-RcA=<L+g38=+
12KYNPWKD^Ye67X:[VKQb1]Y81M_LW<F#_FXCM1M1R9F8NL=,=PH?ZKB-[YY\<Q6
@&S]?f:aGRE<I7YQAIOS9H:^eT/]\>;b.ND;<QVU+W3WI^]Tb;;WU)1TW+>g<,RX
ME6+XR4\c@f[T9X8QIOb9@(72+]I8,M#LgO3a8581K.;F+C29VeaDOd,J,-99EU5
.4[80C4^\8<g58\KG0IE.#GV(6D<38_W)Ia9/K.HbZU>1>@6gIa5)/>:gN_PM1gK
.@-D;M3RCL>8U^3RP2K5<#E^S)aZQg6C?P)3]<6CcU]6M.I]^A9SRbF&,/^Ed&3#
W#aB,c,X&L>.c]dBVBOO54;[a_W(?O?AD/08Hc:HE#,/[UE:22>0O9LZ4L#_2A20
>3J/b(:aV4]K#^cWc-^IbFRQ94[?b:3KPU<bV/L-(U1\7SQKTd-AMaP,Y6/b5?XY
HcN6K0@DaG[^S+MK7AB3F_#,MWg_C81OB_GH2eQ_6HeCKE2gAa+3]Za+W.>0>TER
@M3d?KDG^UI7cO4L80MP)D=8EO7\@UI]#DFbE;ZZ+ZR[b@;(LdUg62F?1?KJKDOL
WNI=<459aJ+_a1EC?P(cIM<b6J];gF_Yf/d>KH=1KgYf063RF(>GR7=L3<>8FE3g
#(<&P=]96<d49[)\-A[0,8QHL2JI^,2<,fdMW-SP3MX+=@O9?5L1;ZSMD/Md+#JR
G2O4.OI?>O8NIJ(#5UMSc#I^[Z2;14S(VY-;<+CUK.+QE[A=FDf:?UAVHB9E(fOP
MBB+K^C(PAN<@O_IDI\=[g-RT_O<4#<;T\&3)<]RAP5[#_0ZS\d\TFHeH6H7g&3&
<>)MZB5)?;KaCATEf5EU]6AAG9#5D\7)dNO:]#KRd;WAQC\HOZLR.H2XWX8WW).2
;RAY1)^0&/UN\4V_A@>WYP/a)B[J/8e-87H+5TcW_)J-3,;-?(36;0ULM6_]gY[@
E\SICL;RLd9D:I<Y8JDM&60g8RUP2.EDdbb4OK9;]dU(KfD?TeMVQ1?JK#B0[JL5
EMaSd8YKaX9F^=H@-M]Z/W?1V:\LK+Z>(Ff4OS55@5]]05ZB/b1?:?>+]7M08#Rd
/<30eSA,F0D5E5]cB3a@?TR])3-^RZLfIB8#50?L]M118,M^VA0JEZgI3MK/.d@8
;,.Z)W_VQC;=-e.TW#2+N&;f=:_3D-UEDa@+MY\6F0KdH<gL+K-MB^8XdBITVBD2
Bb]V;#.1G)UV<ZC7&2QfPKVZCYB>A(Oc45&\EF?XVeCacPIWWfYOGXZBP:-[eH;P
<[B=Z9X&452/VE^=Fc2,4-U8108/dD<ZCGZ:DIC@^X>02@MLFA?G,6_2,7C^AK=4
:74Qd-cA79W.L\9\?N;E7Tc(DTN3UYNV(Ce_>&L8@,E@&=F&F0:AK#dJMf:EBDS8
&#0W03#Kfd)/WF93H[K4d+cS&aeIW-g,B(I?5I5UYAPHM,7#FE(Q(6<HNPI8.Y-g
X=MR:]/UIG\)OC^+QW;b,,DFZeR2[^c]&857YT[/c&I52D)?Fd1]edSU_dCD&&,a
W^:g10g;L0]Fdb/>/bc>dOIN09RGbWAB6=91<4LgR.+ZQJEDQG^NdaWO716(SG07
DIOJ]>Te=-LI@b6.7(E+ZEO=JKYM]U,7#-Z#=0P0V/U9?=^U7Zc<EM(6V8\Z^eb6
[BO:)M\]CSf^9-/.T))E@H[<2QV5=A7JLbFVd1Fc=HTXU=9B;]P?OP7)8f]NVJ_N
Y+W2#;@T5db&Q(Ve(U.,Ne0\7NJ.0J)8]8e8XI@Z3LLfRcab(H:CVRQO(T78a<.#
XCQF8:_P.AVIM/B4.TBV?A?[<P3C^bCecHYVB+2T1436)1^HUc^8g.PZ]^XUTBa<
Q\^+1:LXZ56X??ZZ9IG0+g,Z[1V=gH-]g-5_1+9M.Hb7+-TFe0:_Qc/B\O\,\__.
;GgWd&G+[K1^)3[E(<&BFdT\.83LccXDaEFS2R7GU&1]4IW@V7?daOEY--4B^1<S
d_=U751:b[CK3XUZa[JX-eICQf0^Zed-+-7<EK\HX0bDD;.3H0H-^g+[AdS\LGR)
G\\5R/00;T9(-Aeff4T?&.SS9H-3M\gfLK)_DUHNG,0VTJTF?VKZ(E-Y7LYdZ2=M
=T1)a,c4QVSZGKcV,U>07E9MZ,VaOBH96V4Y0K-^/5R1G8G&@BC8[U(2U:DO2K1N
ZCR=[1VDJP[e;Q1T5GP.dIS\N^MVB&e+(efUbaCNEN73/?#gbJV+EcdJM1d@R=MZ
>G.XG_JNLIZ2>LEM@&23WF.D))Ud:\JEK#-15ZegBJe)IKQ@fQ(]Ud^:<gDKdeP#
TB]ORgQJRHWJ=VX1)]#g^+SBXbR0H+(1eK@3??Dde:RSBZFM<XNbW-&Va/(D=GPF
M?cL1EKD:[WQ>Xd_7[(:QNEYB1EFg)b9QG\TW2>]#(Y9[S_.[E>76H@KZ7)XYdDU
;_JU:W>]Cf<ZS^3]0eSFS,<>;]]Y,Y/Y.MA+F;F0a@#YRDL18_JCe\9-:Y2:2^05
_R^GJ-g+SN+/9R=dA\d^9^SE&.LG9^c]e\ZQ2]MM/[7G2YggaM\#2V9NaD)X\FTX
G+fdG?agb-[T)cUUX)1d^bdV)Pad2>6<WdL?e_[Vc#F_8]LW(b_5-BeKQ[GEX&VT
SL8)26e8@[0aD3TMfY>S>36CAV(5fHZ7>&)HX<+3<1^=&()\#,<W83gJ^3Be(1OA
6ObESJZ[&Y9YYR\NMF\02VfgGTY:_OWI\>S<d>TcK&P)P)2Hd32MNfa^9\I6f2+8
6AJQI6:O?]\<PO9<dFQ<MeD8g3dAOc==f)/\,UUg2WR4@3GG2/<aHd(ST000^)3Z
4IR?<?aDQeWB4cRPD<MDg94RIfP<_0P.2K@gM)=bYb81#A,:;Q#K]B\b8GNeENHX
4)-2H7J+,8PXeEX#A&/E9:W?FWf3e?C##[UL>/V;(B,\.+Ge7PIB\\_W=8Q=PZ>c
_@C_L3K;D((,KZU](L>-NO6T:300,PJ+c4:D[GN/Ndg.7a;\;L=#]U<7dVb3\K3B
XWb>L,^ANTK_5ad;GgWfd-c<==;MgWbN5c_X<H6=V@+__-];;aE:V;Y)=+>1ac,N
K@:(JI5?IE#?43)dM>.JUb55,(Z7:N[]G@FYE.T-Oa<a1a^:-U-\5)KVIe:=95\J
ENP[F(?Y@=5Cd(:D:Y6g5eaM?gaYefR)UY=V9(P-fH^XTI@@>:Jba]8/Aa]?9/V8
+d-@(]GbJ9)g(^CR17ccVE,Lb1KKO>&UQVLCNU:DT]+fe>K)W?>Gf(\O++5e:bHQ
7/O?bTe)8_@3F#3/(&g_+R@.\R_g]J7JY:DR6J/?ZC77X,#T=AW8dXE=:X23Y6/C
Q>AFff=(EC+LMM>PeG>2b1,?_^V5S;N09#22M3AVER22^/KLL(&N,DH50cIEKZ(R
+6=N=@6N;@M&]HRZ?(c\cK/IdM#W#?@)?[^b.G/P]7\:JT&+YX;Qf5MI&CMHX9YG
DGH]_I#GT420#OKaTcUY;fW:PR9(a@H.7#>5;B:,ZW?F-\=)P(39\PAcK0J<E981
YEH[MYZNQ(e^Wd-LTbf+.7UGSX1VZDYb8T:AA&bX>L3?62J\8V;2<dWZXceLYP5d
)Y<I1>b\9MH15C^eW+d>XA)b(f1-a/GV?4,a_ZDO?S<Y4]IHd#]>d_J=<(MM/0IY
G;8V/<0[B#cRB.M]BHK:E3G2B3[fMLZ+R>+=4)D5:c-8Q2+@O#?\40d8\[<[^&>#
G\-3_d7H06^=8Y_>UcJ)IAOVeO>#0=cCPCL&F<bR.>78X2U_6H^?RO0>:YB:W1c0
6]W.-\1bc_IP6TeE)9)\,A&K@17;A0(5SN/?]6?0aJK:YLab0/PR28/HVHG-;X6#
_6=.TbF40EKfO>@<Z:B:>^8+;c50acSg9J7JS:IDD3_0/]^Gf3Z=1Fa1#,_ZG0T<
aD<YfdeF;BA0PX+GYXVZdb6b8R:@(GgNW8[VK^S:bX4ZW+We+-<_?^O#3F4R@AU:
bJ4GMeP>PZ^d.K>3EP3>3fP4Q80TKSVTYa2(.3c,>b;(O>QEVX@Y]-7Fb-Z3c^1S
4W]Xg2V=/>)P1.4Fc6S)BIPJ/HOT9:065CV@@-#99g@RMB<b4DQU+QZg&2ERFM;N
SZ+]dV;?KWc0YXGAL/3XI?S_HWOYE=9@:1Y1FGI6X;TBJG5F;AV\SM7b10_&RVE2
WX]]V2F6;U,J.Q4DT6#cO:R=T^Qe4B3UW8=?1SOQ5.?+.=-&XPT3SO0RK1+>1:28
N2Z##,a4TV(6ae^gc;THZ2[8g4FI7H(c4GgQ:[FWO9QV:QVZ2^JV^XX^#-.Q7?E^
\6#<^V70dRA6POR=-ZXD2cF,X75b0g7DU&g5+Jc4^+#6RF_>67OYg7ER@VGbTW;S
IU3AOe=SO2P9,+=>P26<@,DQC47_cR5OVF>J8QA)D8ULRGHGGW<W8@09)&A6JaL-
W;C^<B)CNb:Ug7#0GM]#1NFKLP<Gd7_Q4?].9W,T@=<bHEH@(X+2K93XC5^f>]>6
G)?MFDG6Y8TH>;2NJ<H[#J?GN/d0>d_[+6dZ++7W86L2^D2-XK0d.T,N=/A@<4Q6
PT12[>a_Dg,&X][bATUd7(CcB^f)8?[?1OXb)+KKW/,\-#;5N&eGY+6IW/5@Q[4K
>(\<;\b-K2M)7gH)>g1A2WN>P8HD79f7gGC^8ELR4BM4DY[YAUER;>(#WA^A/b-V
?BFQ.&^-3Fee#VDMABM#RA1Y9KAQD),(Cd5:T6gQX\S<8U3AMMa<RSH/VIF-TFU,
d>EKdC00W8^W]OY&\RQ>D&9:&VDF9_EO-33+_Y+7_MB(d:T>RC(9[.YMZ9/(AVQb
e>/g[gB2Y)Jcb-N/b9.GQQ:_?Y,Qc?BI?bTR,d,Z.E0FWE>MVLK]DOYc#SYN9&Jg
bODd;+T0T0D\f=T79Q6cGN=Jf]BTNY[EV0LLWN>UKcZbC35\:?VMGU=[-4^<aD>.
MV:55c&+cLCVHL]6-C3M>=NUHZRS7c@F^c0@<MC#.;R:WU+BBb520L2gWQ<MEP&c
I5^QdES2K_2)E3#WD=gYGD4:MZ4Q..4D-U:<00EcYYF4W;Sf)I=S<B>bIP5/C7\:
<Yd[Y+@f07+<DBYPXc[F#YIJ^[(.SM6#XSNK\Z+5^A82cX+36]IOEBGFLfQ(F=OE
JRE;[KD6X&@3TZ][9Qa55<e;IUCdG7.-3NDJ(+BM3QKfV16&WIN);:A.,9^-c_Z>
C--3@RDa./ZE>5Ze1>&\D3,Ub3bgYe0U^(ZH\YL1ZVBL30^<0OK?(JXMHHD]T.8D
V(A&5Rb.^3cC(4g<G/GfZQ?]:Xd_K7_V76b/,+<GS_e)/E#]:=\KOG6DM_SG9U7B
ZPeY^.T&:&fG:RR[M]475R,fX,Z>I6Pb<G3Z+A5.gc_C8MM8_<Vc+J:2d00\[K:)
HeN/gF>UHgOVY6Yce/;@EbgJ.O(,<\,bQ#JMa.&cD@H;5Wc<adD3WKBDOSa^0]SH
YK^b-)>FOE.:d=DAV=SUJ>DYX.Z^[(E,b^@BKH[ABBORN5ET]d5L(1#3N1CN@;43
Z6NC.(C6NMWY/<4P0.GS:,\]V+/7X^AXB@2(Of05<CF-JT/^,A?L:WHOL.@L[1W3
SM:B+<aXKB7^\[#G9:A?gOQ\7=dC)VYg_?^[gKIb7[QF#SbX=/<C+TY(@Q#g5Z0J
eeAJ(_#?SLf\I&TFVI^II(Q]EKQ]+>)UQ,eFLS&.C6J[C&4M^Ua+UEGQ?/.@D.U0
B@=LGLEO7(W+^dI>M=[YAXFXZGKaASI;G:ISg^6]CH[S0QJX;f5817[?A3(K)[XQ
c@>[aYe[2DKR;42Cf^C>a1-]0F)eFPRT0CSW2:?9_bYP<c@2?8?Na;S<2E7F(&^D
V;5#-8&IO4/bCN4W+WJL_KTSg/0Q_1P_V0a7MO,SD1YT/Z96#N8DJ67;MA7JI]?R
XDdP=\A(b5D<D^@^4^+8#f?SZf705C3aO25X5?_:]]+CSO)&+//7+Z>O=aO+dfKg
K.a@3JFHF(\Fd;7JH0C<+eN1\e-+:GE=0KV0LcEXLFX/UVUf2XE:[8>eZ<7@0&-F
NX3L:_&Yb#.N72J^#W=6L?0P(BO=(VC8eO9>(N]/^_SV[G9:3AMF[_4M-Gc0Ada:
3c:T6=C,U)PRKDNJ3<APJ,@1gN=7bg.(JKBH?MJc=M^8Z\1\[?a[XU-T+D>O;3Eg
Mc7WN[+fQPT]R0&GVaGWUdC?KS1]HQP)@632J2JD\U[4)7:H<[^WbK6R+^Y=9_4f
J.E_I48[Q=IP]M@O=H&9g\_O=.<)U?^-/E-9cPe.J;&?DR>[3(+6Ua(:CQ6b[O,J
O./__ReT5W0=ZXX9N:WJ;<f+Bf7cV26RXW#0gA4MPK-#>R[bR1-Td2K@^CRc.\8b
,KV/V[W/?+U\P=S+BN(T5Q3]T+AFMY+:^@?LZA0Qc0WL@e;M4+)GU+[<N@4TT7+&
I1@2-7-8=YYU,B,g@&&Z]#C<I7O_XE4,BOb_X+H9+G6eKJW/\ggSd^@Q9]/b69MA
M@c;\=;aDF6B]AdUJQ8N,JCDI99P2XZ>4JP@\+Q+(1GQ?VAD#,FGC6/fc2L>+]IC
T]-60XKbH3J_BRa0>.<N2Q(6geVf4@V6GE=9GN8B;AbVXb>)gA17#_cZ+-?f6^HD
@AJYZT.&15F29AEMEL\/a4LFL<KQILJ225+]TP:NTY@-b2e//?0S?e8B3C;ME)E5
50M;3@U9PV+O?(3ffJH;J)WX^@4c@/&G<9f,[Ne#OEM&gJ_JF9)UVAHY,<2Oa&aV
86ODHAMZ;1(P<ROEWT+B>CFeED&D#3U>M;dAQbG9a9I74J?]KEWg\8A?f:aFTW,U
M>3KcfN8(385/#aMLcagKMN4-#e,.SW8Z+ECYJXfg(bT/JP6MY1Scc0.f3)V/f\S
?R&(B-1P7=E\VX9=?GD1g/@0H7Ef:Z.=/0#@3\:b.T)@8,71YH@UC0Hd<g#O.O5?
>2U=bHNX3^e9MLKbLaG##ZHTg2U[Yd6P^a=7e[Nf8e<FSHXL:_++bN.f;ID\B1.C
>EaER9b5:M[IZSP7fLfO-PZ;OOSS3#M[bBHZ;-AUZC8)3K8T2S6ZAG?b[&d5\B7,
ER\d2LG;=A_B6S2:WE)RLN)b@7QG_-L;U/88FAdXZ>RdV1#4DY+4(:2AR_WZ3Wd1
(R2If/a^,0Ke>)F3[LS_?5=MfZG&4Y#<=YKKVK:(5[)X[gcdf+E1VS3E6D<Ed9N6
^\(<&cDS1Q29<\37+BVf@Z=_A4UU2[#Fd]G[-:aE)RJW&]Wc1,=I?/ad5cb.XOG@
/gYH#?@V[&Z2V<N(_HP&;8g>V[ZT+VF4JM[UV^7U([d4,4GV[DM.W+]<c]R5>Q_K
]D5CH79_<Q4f2^4:MefVc+\PQ8C)0(/G>=C.fbIDg_^H=Cca.eT61)<MKGaA8/?/
-T?3S)TU&<.NH1NYbZ[A#A;^HfTT.cGBS1#BgXZ[]E7_RG>ZWCD\aA.HF?^9?A0_
G.BMg=W)CXJ)+V;?RIB6EW+4JL8(FX5C3XfXE(=D_)TN5bGdS)eBPKLZR<=NfGE]
P_2]R:CLOCXg)V2,S6RDO+OA.c=M<)QIPQ7@M)6aVdHP9cE)&[9XRE179V11B9N8
CSO.:9?M-_QY;(_+CVdJDN;^a<cV\_O0-QLK[M1)Mb=<5VK\DW;8<^g1@6Md^A2,
9>H8YHfPQ\Naf<T#^&P@9W2gU2P7E)aXY/:_\O)CBANDBfHa4,-f.W_(\.]V,<EF
^3_COBH\II#SD2-@.(YIB;3HO134A,[G6;:=/_GT^cQ\U>60X99\#?I82WI3DFW_
BA;I?aV073/3-/S740GYMG+<Q.WB;PbXdg<Bf8YJ3D4/.eFNdH/TA<5RSa:<EZ=.
IR.Xe);DWRg;HIee@=444:d-OXLV7F3aVYW=NPPNc6.)DDa+C9E7^XOWTSe)E8g;
cDW?5M>aGB@K0++ZIg5G<WNQ6DDOOcS90T6Q@[/1L.&56BEH0c6?J[]VL-+9]/=Z
&6&:\-+^;a0YM9XJ5#839-/EX#g21#J7Z2>4W0</,2eI-EAS8fWES^_)[U,A@UOX
R0ePNLJY?f)R2MaeO>V>;N#B1<D.U9AZ4CFT-SE7da/F^5)UY(=2/XM<;fb<6</^
0-S4_1/O?;Df5JODUV?L-7aRR-N1>6KV0DO<f#&NDSJYHV1Q#X77A09S99VNQ2B+
S=#X--B3;U=a26&)c\T,0I_7.__J<=W(YQ:A6<J>LTcG_L<H?15.b9)f&6C/A]K(
&&1T/21&g\K?>+#U>XaeKeE1J;UZU-S2=ZBC,)^Qf#G,daKCDY4\Z1.XdQ\<9+4G
TcQdV?d4&YO7E[3S2YJ;8S(];VC2CZ5]EOW0T&(>D,Z(6NV&HM;fTOAU=D-S14Z<
9c\;Ya>JT+W#XOE<_U,JfOLM2+GDE_N[;CXR3_/2M@+OZH4AXG:X:P_+]:Ae&FX@
@^f7:.Z.bDGEXeG.6/R_Le:YT]ff?L5V[]K?=,_eEE;X5.&VYDWY7c.P/ZP\AR1P
OB8We5W@6a_;c/HN9^[d3,DbW/KF&\FP@M(U_<9987&EfIG+V;-]aO6GMQ6QI0,@
bAHT3=6#YaA[4N)@)2)4W75-PJ:#SSd1OM+3YQHGL<&Q9H.30=g1S59PTfgVM=N9
/EYb7HJKISf,YG\D0X>Je937R^LX-@B9c&E:gJUd[KJN(-#TO+NZ>:]fWKZLTA^1
5_c-bJUHOB<T3=;Q#25MSA)LHV>Dea]FX82/2T(P6HIE/]d1]@e;aUfBd6HI-:dW
Y&a3)gR?AgVE\GX<#K&.<S5KM#YE@2@]4PQf]WN<R+a6+AfT/;82SUW6XQdC_/Ad
.+)FB+QGRZDU3SfSVNeYfG_6a9GaDW\[DR;CRJ/NB8FcZ)U5JV4L0(IZ/Gd#cb?E
2<1#^DeGUbR+Q^ICJH9#N+3C/KA>Ed<VA+I)7L<.f3NKAG;Q)ANWgeBTJ2fREc?W
Q8,G:W<a.,I:OK6>cYFV8JO1[V7C]cMd?U]0Z77:cB-#<24dV;0;QYLb;;Z].R><
YC54b=/M[P_&WKG6?d?\/_:^?cdH4<LFO\64@4S\WIJ(Wg1^c4]N/[31LX)aMBe^
0U:6WcbAca]Ld-LLaSXE]WS7^&f)VBHf,>#5SLeBZTRD-SG\S=>6258OY80X>PN/
-8:+S@91b.#1K/OIa^3.PPeRP>UH+g[2TYZ>;+cDI9[YAZ+fce>E.B9R\6#a0=^Y
1e(23OW>:6@eXL26Z;c-:]4;K0IIKg2^8HR8:;W.PB@(^R<M59[UUgAI@e.0Gcg3
CWa,)/J3B93f1I]9:g3QF-e9=+ED6Gg:XFLL]];NCMZT^eNR[WL0<[6Uae?g6dW7
K(J.=7.G+RMG24\A@DY:]ZP^f8Mg[514G87/g\ec^7dSNbW2SQRD:5N[J,E/-3O9
:-e(@9<P>K[5YTD1>P,D@=\T#P,<>N9.beQ]>fSNb\IF_6dCD:S2)FgW&ZL2FQOC
)@+ATV4CS5S&b9L\0Y+UN>&.N.I+O:1XWc,G[[5g>GUKICYK<O8Sg1+]WRL;2F]\
6915Yd6N1]D55MGV?Kf4NA2?^2[=Ed/&#(c>EQ#-;.fHVYZ_L3Nd\M?O_945c1<9
.V5S<>UN_Je.F(]J8_R)L2S+bR\c]7UBQE8U^a3cYJ)I.01f[eK^]3,3d]A#=L]2
^b4FfL?eZD_/EdYO[XOX]&,?Vd2D2Z;3D<OKF:D6^b2LP\]@&;]efX;fPgD:cKN(
(4?.PeECC.)c#<6(A?FPWIWFTbTR+5(SegQ]D31[J\1(/@.XDJ52_HV5DP2V3[Wa
_c8JH=0L>SIYNXfU:1GUT2>4P6PEbJJ/>[_Q:P0MI[?\J>6-8R^D&1[#KUCc4OEb
87XO-1E9.J&))2Nf+O1g1RXXEIS6TdY42cg.A;1+2W6<BSg9CN_/-]a@@DEK:b&g
R4X9A5R<U3af1de#X_^@C@E0NXe_JSc^&=dJMDA;Z1H2WKEfH?N1#N/CU[e-:C4_
ILbIC&U6bfH)\\efd>O/3RSS1XWAZE11eQeBRQRC^Q\VbC4X8E^<->URbf\P3S2#
..I_\M)8VMG&F)IKI_8=,9MKGYS1fL5(A+CfJ_OW&:KN5,E37_-1.@3<[3EJ7Ad?
e/;18IT+4C@ZSbR4a2cXZ^)@34J,0=&[U(-.YeaS_;P45@U6YX<7@Tb[>Qf7<4c:
+@0#Y=:<?<Z/75Q3348SN]R&+S.aCA\a<Y95-/F1STT),L=O2,;,+J[CI&dVJ?<)
TSL:K5,-WXY1/bUFM8LcVJ]0F64A[6BcHSAYc6Q+aSf>:R5QH>?G=+02I6ZVRfV#
NfP4?A8FN^N>Q<8a5gX<U663cTd>)6J/4g6I?P8@&)25g<X,L5SA\UW_@/],=<\:
Jb1P8L8TdgK,,W?2E]>O8HPAL/(g4I1B[.=&DgM=X3f[C)+e&MDF.UOM^Q3@?X\M
VY@FU5Lc8eRM/7D][4Seg)[EZ)Y8,@OO_W(<c2c)UgV27/IUR:\-#@#]PMNVNb0O
d?X\4<?TDCLB3O&?eY#86OEWA<(ALS#)12FXTXC;d-Dc[:@CDZFD4UO=DGV@JJRB
5I)/,>+(=f9^HKYBU3Tff58OTf8AUfONO>debLE.8.3_f=Q=L16\5+KFTg>IbS0G
9Q5(1SNd(OCEVL>+1474#TSCZe#N4AH@/H/9b;Q_1T+U;UaT5gf:Z5)[fON_bB+7
S6.X.@J2@=O;ZZS.?VDOfc&5gJS\^N(M-DeO6IfXZV=b(74:Z[Zb?;;[BG]II>X9
&db-aTR#\>O3#EfKJB;OdTU64G+eHbK2]RQ6=?\K,[A@IQ2J?5N]5+Se>A[?VZ](
YE:[17OBP?5J()VAgX+@ONa0e;M,:Y7@V_VAdgf9EAB7NK<UggTe9V@SV_(5gMD7
E\BS7V_Q-YO8,I_DS#Q._6<@d,L17,fIC-01_PQ)>ef<5H9RJ-C&S:--=Y#Wb/Xc
NZKSEZ(IE><Y8Vf3,WOO=RaGc\63K.HeH(XDX7)K8IWH8X2cVS?+J,V\NYYMTVPS
47Rg9FNO:0(I8S-QPWY1>F9F4_PIRYXa6;eM4.UN/9WH]J]V:.+b9>?0MH9]X0>Y
;N6OA7,I,HLcJ^\;8](JD&#C.CO^R(7,A.]CWTfO]^ONP1K-L?)->T@3:;<[bMc3
@,]0YL9b<6FI:IfScQ:0.]]MI<XBFd2DR;WWMO#KDL=;:L7Og\QGP(8\AbUYI3@B
3g0-A05]NK:/<<F1a8NOL<Z>ISQ^-SZSFWDIe.35V^/MeKa3O0cZ]37,dVU:<RJf
9UX672?\(8[@PaZ<8A+2H>X?dX4KEAD))B2,WD;8)U_b(KQOdcD<9cF3<-fXO.\S
&B20GG#&0/AW12G?@a2QD7-\RLP@86Q:aHDLY,5#eacBZ^^N60<O0?SQEF=2YQ_D
R3e8Ofa]>]6EO:IK2DO35]cKg2TVWO8]Ya3[H4B)PN<E^RCJV^\1NbU#.6^.&ZHZ
cgYKT9DGgH#/d.X-g?U=,gP+4@5\LFP47g/-8JPPOBL0S2&FfHQ<B]<+;WCYAcK&
J-AH/YYDKCV:S9W^B3&S<;EP-)HILT862F=O(B+=S4dfTL0Tg2/C19[9-U?(^R(3
Dd5O+J:]7M(Z.[J)E0ZS)XPA9981\#J)FdfS@^K03.?\+PL+]24P=-9)<OJTe]=0
>LbFUE@Rb:8(bM@4_WA)-5d:aB#F8V[P,<_2fg:=K-N_LYM\F48O@&>^=?#\\L)^
V4LFU@-aQgD?H<g.B+?/.P2-NL?9L.Lb,GNgF<4J3ZAN[8.bS-[82(=R=V7@Ugg3
?KDOZ^]]U,dUS?J6C)bWfe(=8XN#Q&<0H7W&\G2_@5Z,PAL_B249]/@A43PO(dPT
^cWLBd-?J&PK[FbPQ#QG^IK.>VB<QS];5C5e;2,\0Y_bR-.Nf4+e5?/8O]L]>IeD
]#,^KETd6I(MI;Q/;V)FO,\e[27OeGeU@b;aS<A<HZX.#(TL/SW\dYEYWNOV]L3-
=(c,0MA<0da?gIX:TZF@3+&e?2+fdLQWdO;QSB8+c2M/<5F8G,VX^N1a])c5F&c?
),b1]2:I;cg+Q5T4<6f7(J3^]C&f1T.e/4aH>G]\]d.0JI_K\]X/[K[<6<61KR\/
Y&L_gQH/OTPEQ;I)AU,:@D2;^5M;_CBB8C6Tge\M\S?ZX8fBeOK0&EDM(KMgD#cT
\.+S;C8@YZNEC,M-SdSdRF+K51^).9[5?;TA1M]--&=KNQ::E2.S]6FB/aY\@&F=
)(<Pc/H,@#UA17T:Q7\bZZ3>[;26P)KLI[8@,-dN:c?e>P[8CE?@f3)F2I<a8+e\
Bg(eEUZ4(&-(8Z4W..[CM]-/=bS7f6->L8?=B=LR6GZ@-YO6(B;c;VPWC4eN70K8
?dH^:dc,5U)Q:KO9:^=E;?=4T:cd68S46_c.aU4a=N1&R\:[1I,)7/aOTZ/QaG-L
]_fPT=+F@[/S)JNTPa?#&>5ReJ&#gGcZP.-(JEEL[[Z(900Ndg>_0gdc&-]#^BUc
;1QcaS3c5e0U:924Tf_5]-a(&M\6<I0_g39#3fA8=/5U]3:fUe3X[P;XM#Q=-.M6
QW,?S8.F91&&/USO>dJ/@Yd?<+BUe]3BAgLA9E+CE.:bIce(I9eEVFLT002\KD@f
DgBI?N(4PB:/dR:O?Y7<JLb?LXECE1J>;#<(GAePJ9GNe8AH3cY&52gNU0FP#DPT
Vcf@N1Q6:>HV9/KH23T=APC\FTJdd559.A?/)Z-H2#N236YE@[geFDS@-JcfYRL/
9\R6O:IBZ4A?=.BO5X<\4IK8I+AObPO1d[H]-@UAfNdQ7TaG#Sd(AdFGY;T)(aS&
XY+7O?UbGMJ_(Y4K<cPH:.&YO(U?8@MBU@PgA?JUX,T^5V5<^G\_TRCg<HR6M)V[
V0ZbIIK<gBA02TNKZSUV?[_9<.]EK&G/4,;V&bG<3YB77QQV9H5\\G_^I572Rb(;
@b:e]7bK-X[eObIE&>M_4XJcbf\/:G2I+?B8;+U8MZ:79_2SK/F<HRH05A98f]L<
eVTU4RV)V>W[183HO.CR\4f2L)[<RO]1a@[56R^eUX[Q]6R@GCXV59Vd]R<^614-
g[1_(U^YZ9L6J_N4,>RC>7gV9)X7LF=2Bc_O?U)g/Sc6ECK>/DOD-/eJ[/7^5^@0
XX#Q/:LO/]e?a=^;Z,=]eBB>e?.-DJ:^eY>_a3g2ZZ<BJGbZ[LJB-F[1b,VPg9?1
FB8:8G?)=SSNbF,R_9B;0?XQWTUXQ=^3@)S62eF9WGGZ.fLZEV^VNWWZ-P3,ZSH;
50>XSO_[KHQbAeMHOBZ.Y,[/44F7F^<0HZZ=W]34,99Dd:YD9dKc>4[-50EEc<^D
a63B,N^_YDXY,fa6:\fJf9(#cSHT2]YJc5]9bH2.e=LV:)AY?.O+Ka(_8:AO(#F[
7TBaUSD^K^P<T&D,VC5U/8c3=Y<Ya,XM#5OIE3N0ZV+?K1,A9#NCVXRSg7@JR39a
;#LK_/Va&/.b3S>9DI(+8N+L#UKd/_R>L;)MJ=W)RR=TS(1aW[_9=fCFd]@5MX;_
P7g_PR8?e-0_K_=\C=3<(1/)&1=G]@^>K;\@C)aA6)]M98R)5=[X2J_5GQ7aC),L
BHXAW)M\a8UbHX-KH:6A-K#?7E30;,(W/3b=.UHZ(\[N8#\N;fIA^fCU2CL85GY&
/XYBE:5:#MCW+Rg/XK(]G&g=_)&+H(6QdPH@E>YW.&a6=(d5=;L-;P-c^SGIIeaT
CMc:[29G1F;gJ&PP0;S6SK]NWJ74V=3LK]:G&a[cU^J81O99,g>-LM72HV22DW/>
+EN:HdQYfM\)g4a@?:V:9/A39(-:+OL:5Z)O<eIa8:B1W[LIE]1E75]#X57LU6C6
1X/OK<\@#@e460&S9/]#WJV8PJ:FRc8ZPCQYN?Ld.0YC-\6La+cb9\(X<BF<>]U5
+bATG@+a4IV+IPXcZ6A_JK7dbbXW-6;dcKa<7<5IQ5SA5>L,OS19N4gbD5]0Q.ZA
fOV#a[J@?\\Da\?C,S_DR-#HY71J9U,2d7_+RF2?=/e4\&7D9V-:_W=_76Taa0R?
&U6XS4BcBG;&C?P#;,G3(f0fK<E,VCf&QO5&\II1(=HK1>/?\:+ZU@afE]ON/D#f
?&81H^T48bX6bP@Y@f+)30RCO0INST./LTHYA9O]a0N#>.=5([aI)RZFWZ&/gI+B
L=#6b\TZO7bAXaB8dO@(b>43A/-_C\01dB2P.[E&>a2aYRG)N3SO5;T&B@b;RaZe
c=R^OXDFM&<O7YXWQQ#96<[AYBN-]>2^C3;/f6J6NX(c+IYSZ\KgAUO).H8]DTdD
OY^f[#a:F=7XLc\[1]1>V>NVOf)VH=-bVfDA+PUU43Q2NN=VQe1^9[M]+<ScaT+<
F3\_;S/CUQHe]7-6(J:HTP,W_;@8^,\5b^-ADbbd2AF0gVN<+&9B)R9#,)REQO,_
6BL=F1B9g<1d5W:IbR_VELOX9-?ec5]5b6;UCL3-_beC4SDU44Z<[U;1G[3eHRa,
gGWBSeeZG\IVQa<_5^T=Ra@B.:D16[aT7^8>>gV\D8WQ5;EQe:XeNW#MF09S@BAc
XY0;16T7EX2NFPCWY>g=#=?T]L;S+RO6d5.f:>#O4[YJ#W6/X/E@gCKD#M1BW@F7
7:OH@UD2Lfg)c1V9E;N\5D]?RI,\d.Q\YO@J21_JJVOUG6Oa]aBVN,GIATH3(gXE
FU=c:E(2S2X96;[?2K0><_L0+LgBG\S;T5Xa6a#MQ3>.I,We5UO<8O/M_dKZBN23
5)SQJKD.2?4TL>@+R#\:\A^2XJ#NLCR;&2IYCg(3fI0Xga.Y6T&+F.PgT9W[#B,)
aW56+)#OH(cPR&KO<>B3UgaW7@O^OT+8G&H(aDaYZ>2C<_TG:8?YS+H.gbHYK38.
VS&(F.[S@2X^S7J>-Ef^T[Y.<<]ZOBAHGC_G&aUFL[WTg4L4(UM0@20DZ+[1F\g;
aYJ>:Vf7JcN]EBU-S1S@V0PI1MQ@PdL50KJJ?MFU]=MBQF_+HP(KfDb:QL\,[A:5
=KfV03M+-;Ie>,^WE4ABOf#g:2D->.3eXL.I))/ZOd1#N3N]?Y8NX^=TSX;<+N:D
;d/@(=9bJAU]Q\aX&_922#&N(;Z[PB1J&Q?@S9)O&]J\6RL(f2>gN)[R)F:.9EXU
g]N&D5)fLE-/ZL4UB1<4AFBQ?O^/WSe]L/KVEYM:W5OKM-1PeH\#/GOS@3MF<\CC
P3-H,N<V+-Z+aOK4L1]2=D-Ng#d0AS69O(2-IOUPB\YY-(8_LRD3N]#(J,g((=>]
[J2gK^2NRK<]+J&S-Y\JI63/cdJ0<4(2]9^S:/8/9Gc-G3W,dWgP?FGf2CK/dd21
9eK9=A./Qf:5e_)FJR@J7T[HB32>c5Q[:5E6?aJec._@\IFeEG@(NQQ6[J[>)PAA
;,ec#^I^N9]9\D>@gX0Y)&::YRDgD&M>=HGIU=U-;>bQ-d92NB_Y7f]6MY/09/Te
>HbaBE9^,9)1ZT^UL2e<OPCFC&IaT5SH>G)L#GNV>,b9CO;Q,/(0AKCa>d_,3gYW
9#F;2Q9D=<.dQBF28d7#(EJB&0P@_BE?Dg79Y(g5UOgS43gcW#^;V\/HO<C8]0eZ
S?6fQ[^N-bWG29bE@[V0gQd#U=2+#8CN4.U,(W7cC:)6,QO(&DeVMD6)B_=<\b9)
].<PgRUIgW3ac?ZV?V@9-&ebP&89fPG+:@&8F.Qdaa?fEF[LHdV_;WU2\\&>K]S9
7>Z=aZ/3P8a[cA&@H.&O)/07<gB<@X8[)06>;S&W<[+T2_B8JNW^:a84VND9,9_&
^JG62_U:Z6,2+^@2=Idc9^RgK6_S.6^HD;@\<J#gI^.Bgc^=^[O(?@H>[Q&3L>-.
5eW[,L&RP,I6>O/QZ<?Kfb3a+I=K20](8NG3Ac,XcUNXJ#4YWb21cSM=/BNB#]M@
-HMK@<GUS@Dd4D[D4,PfMUS,CgPc:@W)8MBI(J4,=5/NJ23J8#Pb\5+M=LYgQgLT
3f;CY?AA7QfAF\3:U/\[],;1-b0AQ<]6U=1IBVcH)9ASQAKGMWR-MZ6(T7)LXGa;
[,\HFA+IgJP.2Ic.9>Q&NbH74N>WRe-/#9?=5d_L>\)?/dCHY(2EW]?]+\L[,=dJ
^O.F@H=+BR[<4GLCN>^UWM<S]Y-QN#=9^GNc/Z/QTe]d(QVYW^3Ic+ZSDK/9;[(<
gW3/8H3Rce0W3=6H[NcG\+]^XP=g2^:4ZJJa<<?KZU7?4@-2#A;,>Z]?4gZ\^f35
981NgTf,&OLZTUW(S+19AfYZR^M<?f_>[/6>+<).gUC0UM==\fTWXB(PBHNPQ=V=
eDJB,^B1b4dC5P-b6MYNXJD9GE=0aSF/gLHDB2<7A68&=cI5gU;9ZE)VIY5aRaPR
+4NQ+c.dgZLT2Id:e\6>FM;3ZIA3a_fDLF:8&5I<@E#aCg:EZ]d\]>aQKM/JNA,d
HbUPTXUK/@C&DX#SVa.LUGg;bFaG11[,;?.>FCIeMW7<^Je.G[+d=ZINA41M,_B9
+N>ER+3=^8eQ1cSaA0GfT-.RS[aE3=U4>B4H&VJ>Y,[ba]EdL\S2cP@.gcTa(IF(
^M^HA&\dYdC7-6>AE_[Kg6N_dc9ba#JAJU/a^CKO,[89WYVRAC68=IPD#a+/#(R;
Q=P<GC[bJ&R,Me8;5(^MdWO)eR;2LdC5=X0?P<@8g/)Dg?;@-Zb5HZSC=0;7A:&#
@@eF]1^0eAKO9N6?U,0?8D1SN9L#RQ,#0])GG2@H_RbXI0BVYLOS(NAVg^MFNL92
EffQ5=NPW8927\,Q+d8K5cW3YfGX?AN?-JbE+F^PBZ>I\MZ^>(Nf(^9RFDL0B3NC
YL5PCcd\d?Y@7CYTORI5a=Be4eVT-?)PfU=#(b3U_1.]7]:]1FX3YG+VMFZ3J116
WZ+#_2,_#R8d8GUPQH7IeJ:cMc,\801?;S7\W[#Pe(dg-+#;ZB+B+<[=H;OF&:8G
MQ;#P>.Wcbc<OXJ+AS,.2W]4bLc-R+bg-NCg#&)88UQ16J[M-P\RaH@/11#CeUWK
H2<MJ;=ENC>SgQV_I>I(ag6,D.cBYUL,,VU7KJN:&2N_>;d/BYORK6]JE.g^^R0Y
0e\K^GYAH6OY:c2C.:\a8)#+KH54>IY@SVf+ZXO]I.ZcHU]Y[K@^]O35B7c3U](N
70#b(\+YL==H,g@I788)TaPXJU_6;DBVOF;M4WELYPf#L_4BEK^fM7T4cU;-;#[a
BS[@Ue&C#M@&@;d&^)7]JOIePN51#d^33a+ZP5KffH<)D-cF]BMF?A)A51N>.B3/
NA+JYJ595<XY_YB^^(gRX_8#]0]&=]J20S\RD5[1X@f@N2fb_JBP]N7U@]/:c<QS
NC1fS(,7KY&];HBc]Q7SP;+2[4P@0-KF;f9fD<.PF/gY+@8Gb#<R]2c^HHJb]5C=
,KNc+QFDZ[HgJZY@_TH(_9CU_.U@M?1.EI2&I7G6>1-GI4cG,Z,(/;HE5I0EZZKD
MCNNT)gI/9]f4SI2a8^,S_^6KYPLU/(\Rd)_-#f<YIH:8UT7.WOb=gS\eV,5?4Lc
3_e->+IW/c9_F,P(<)DK1a9^24),gF_b6,.8N6;3gA6(((0_g2S:(.V3INL=.V^@
@\5\dUOb7P]&W#EK^@R]:VgKX+a(QCF@HgR=4d\aF=AFIW5#-A.85A?KgL#??PX/
7KA:G<;U?c.L(Rf<CI;LPbE2B#V(;YbDG-D=)eT2DZH;aU\#/1:_\e2MJ]1=R>_,
-4?[_JCCc.Z<\9O4PF7[b#K1(K.1d2#1.(..[QBYU6U>[D))_bEg#c.2_dY>+[-H
0C1:Z(?&3SfLK6,bdNW2H=+E9;gGU<ag5=RZe=7R>,+KL=7TR[)&T(1d.\)LdUNU
ZZ?F#]a9ET[F)V7@XBN7ZOL7Fb&O7/-756TOE3edGD[7#:\&JB/R(+(0])2V>T56
@D<b=I-0YN=A3eS/.<:)Hf=4&ZEQG8(aW@cO3GPQX3?(WVcL,V?GdDFTf09&0KAA
MENID^&GLRT1/ZV7[_&M_(12BE3IQ[gbZAO=70:&UH(BOO[c=aIfT&JYN>dST0[S
HC6FV>dU?)NedX3;.<46T,J@SF8B4IX;G4?958EZ.;32fQA).?>Q;&E4&.cKUM#A
+;MR.?ZUD^KDD7#8/cMWaKX:b&7d5KA0(g6?4@?g]0-^;QE\GRg&D6SL62?cG.g_
&,ZX8KCbF0GfUg\[2KaL9,0VGOd([=S48]GYEA8=<X^G4eJcgVYBCH+cMCe<.A+?
WKb-N#D]1E3)cIHC.V?I]_7^^PW91DTFcSZA5+QY4/#,Ie<X[,d\<;bH@629b=5,
0D[1dR/M)Q5[QAb7c.JFG5f/fFTZQ7,dV1J0I@cIa/;BI7+?\78N\g]VAPD.7,4:
/9A1Kc<M&O#>5dU,NCL+ebTETB(9/e?)?>+\3cP;0K?C6Ub^c=GONF:0=_^[,/0B
,AEB6f/3f1\,61UC0CKaNRKDB5W3Lf)T(P#K-XSd(D]U76CQJaLZ2SW\B(OCf>Uf
7CRAF&Md[73cIU-=)8f86PN1GJ/S4?)9D3fX2b;=<@T2ceF2d:\L;d#-NH12S)<#
#I2:MWQBXecF0V@H.9&ebFV#SD+e.ZF8;:gVY-VTA>,3B?3\U,(0,TL4^fU0_\[_
]FCeH?/91FLg\]M&N@=^&+\cf@0U.Nf/5WA7WB/A=@Z#L,5F(5HS])?Z58c#7=B_
\:E7/EGD?1Q8GFa4:@:?.GBW<cAJ1f8?1?QR5-.RZ,UX7L((<Jf53NaC5SN1._R_
P7PWb?L=FU-A,,La,/V^6T_7A(1?dWcaN8NZf,03(6DWgV/I[0b2D9GVdXN=VZ^Z
2V0GdH87]/BDOU@#<KBKVQXFANg+O^[,3RN+8083@X>:Zg5SR)GTM;J)2S]>XN(U
=EXG:DQ2O8:#P5P^.121N,bY(CV=,0\_G4ZQFREBG4.@]J9@FM_@?IQfEPf]]]N3
&6)9Uc]01NAV7P[@91EU:OX[B=fBbLaOOAMIVae;CXdMg_TS+R.WCMEAI_[[4g@-
410/UW^MN^d;.F+^9NG(5:48P]8a_PLWA//c:XD/16B.N&Mb8EIM9^S7C-RI]=/A
+?2&1LKM_f@>@>EA,+g^?=1eFM(AP_NJEH#XT+J<&a#/(&7N6J:L_LJA]M2Y-cL[
g-;.b.8V75/FfbOY+G_8)10bLLA,VEg9\;I.OR^/;?F?FTB42Rd5F#[(/JUXOK)a
6AA<R.Xb@@/;D[,7_8N[g./I7RVGAS=4_XHOA,:1F,H/3Rgf8B?Y#J.<1U2,/I<f
N&e4Rf)aB:6HdA_ef3/&ZK5V)\b/&RN?8CEVPe9@([@B8N&ZRVDMD,M:LfX:\^GO
[5/Vfca6[UY+]N7FMSdbLS1ge4UW6I4V:(fS]9D.JW1R:(J9VYF,)6a_@W\GA:TK
H<K30bfC2aEFV-M;3=6)59Q(1?.,GO+PBB\>SMg?W6Zb_+MIfC@(#YVVY.?;I-P.
g@(b]-Y?.[X9H7]bc,BF4[+RAe?05;a<gLVW.VF1f?AS/g\15S-f/GMW0LXTH-^)
f^bbRP5?cTW;C6SX3<.LW8;+-bT4=P;A27WcP&?EX_S35WP2QE-Pd\W;0+:()^@+
_YYV&VAfHFRVV2U<,\V?Sd;aQA:B;MAU3#a6=[0(WR#+AZb6g6K-d2b?##bRYAA=
af_QCR@[MCcd6OgcP(=HW2^/Jc4J)D)N,gbJF9[-(CX<cEH9TAL.K\>X-1d@MbZU
1X@DgBAD]U&M[4=6?)/X0@1&EKX&TU8A5cEY:Q5&0)-,S^W9fZS:XUA=d=N@?eKQ
JF3KI))+F-R^WfH1g?+3JaeCXAS6WP9?FD[<Zd>7JO.U]?/DC2E/g+XKa)@I.G&c
7L=T\EF<(^2LL57.UL][H+4bU7N,c&RW4=5581=N.Na?8I+G7A8Q+TLbb&Z4f=X+
V>)a?X+/A6;2VM[O(1#<T;FLX\EC-1<PGdc<7];6[]>UD8(:(;[]MDV44bAF;FD&
g1CB4GYFd=GR.N(S+19(PcF\5BXNPG[T5&<^dBOE:,H.4@:d7?TO0Qg/Q9W,V=_+
7QT8)R7ZHb?S_X?FZ/UX<?.B_EA=Je>EJ(14(0f]EWY2Q[7QTZe^f.XJ>JSQV_37
:_0O?b08QdR&B;(cbdBR/#U=_]DMAT57-1+0_UCWc(.a[)5F]d(N;g)DCEF)e+GG
1Z,e1MC\QOC2,[UYHZ==ZOF8RKF41UPV7De1\6O_=C?fQd-gPZTW\g]DK8TE>/#a
FB,)]:NZ]VUC^dWNc_B(]5bVH>c@\g#FT9&>@S=70NXVbZ(O)EB_KL#9(1AfeeY[
RQZB;;J8UD^U7(8G&9.?40CM9;.];17g>^6f7XJf:<YT^6V/42)MS,gIITWA)I?L
HP;S1.BGJ20:\QK]9B-5]F46ASBV?6HO66LXXEfM+H5a]=,5UU:Zca^--70DeK&3
0N+^aRTCYQaC>b6RPa\-:RE^c=/FZSeP^V>B+IPOAb(#,>JY^^a+?5];P47L)f@]
77UQV^EZ^YA+W][:_Z63#3PgF@^ISfN;HXfHR>M8EF2EW,7CS^]cJP93]PLXF>>d
-TC4[8A73e45G6W6A,bE<@,Y.[>J_,9YL]H3-@JB+\L#@C&<:B11RDX:bDI+/e#b
@R?9:f84_#g5HYQR]T)a(E-LeEM23VB[#:F=>SC@AfN33YOL5.Z9b4MKE[&7Kfe/
E,0[IV2M2X(NeET[Xe5-[-QX.75XI5_bG36X=^bO_[6ABW/]?DTY&dS07-PdIK,P
J@ZX:^#=X</AWH7WEJW4Z)K=X2X2MJZWE1&B0VN6KW.H;@Z9PLLQ.3TV/g#E>c/5
6Q.RVB^?SR&>_X>^KX[YM237^GK21=J/4?EcGS3OD1/e0G<7@=d1)GM[8A&bY401
0dP&C&a@G9#,H:HK:93b+<@&3&3]a-3WH<XY/ZWK?7KA]5RFQSI0P7&g#dBS)V;&
U709&\7AG=BCQ,)J3.A?.KXFHU#ELV8O31(S7Y0@S<B/-CD2+D/<<-,NAfY:2dL?
9d=8[&Na.3:9II/#___)bMb2P8_c-b8d,O)24\>eU>RLf##:8J=GE)^./=JP/M:R
fb(K(](XYG:BIXUB+-[C^#eZ8^:N@g779::&eA6>QN>XNW?I=<,Ceb31,D_OgS&&
MbS=JeKgV.QOcN=Q;IK6.@b^QN#b2&88&KAOe<IfQc58;#N2G=M43B.6<+:-&U:Z
5Uc3_0OZ&cfZYTW<P<@GHV(#8J;Q>#e<)e9RZ.==W9JL.?M0^9(W=ZV63FIH<2MI
A]YL:YUBS^PP:fI]3N_OdbJaR0V,Db7CV._B>3d,2[U&7S1E&c/C5/HH,IDe#\#1
DK?D?XK#3^)[ee))@S&<6XN)B)4&FBeE\:=3Ab84(.a:=UT^E&MGT1Z/@&I1=(7O
7&BMA^c(=>5U:#aE-7@^EI1:]XV##@5.#.RQK_5O;U7ZE:S5-C73=3GQ-P+>59,W
[9e/aNEF&A3a2ZN,^IbQL:DXF(PA58OB9I7TEQ1dQ0^<7QRQ<CZ4=VQb=c^R^Y?S
N95[Z.]S?/d344/+IN=J>-.(W^N)/Te[OWSQ=NYPTO6KCWaQHV4#,4D?@5VeU@@G
ABE_PS/DBO^\KdAWQ-6E5(T,^ZFM2<O7TZ8@T/.0O<UE+;cMbV0R,K71:0JN9Z8#
Of7GOgb=ZP?g=7\I2e0Y.b2Dd8d2>>ZY7WP8W3KPT9S1^VRM6X+(9N,R;5e5S+?e
7_,8Z_,AG:bD]JCPgY_11Z=YX;:&[EE9[>fUVHd\7/HR@MZ9.MHP5;_?)IWLL;HZ
_QUU_9-FPU?aW-J(OaL,7^ga?eK-28+O-;_N,4Z(>G[VaDa(6>cJOXPc(T,#W58)
CE(b3;R>B;D>9?_B\T4M8P8EcAB6&5UKM1\H?7-;^K^-2I@,\F2+NTB>Q&3(4]<R
^B67G9<VKc#<9HA_C#^P:f3e@FM224<?FX&)YN?<)GV2@,bRJ4EZ/,Z::+\QdZPV
e.<gS1aOg6NY@=-PPT--YQB\,KbTRGRN]0cNZ_a@SCgc9;_+4K#gR-J^#dK_+G]S
>1H#8e1S4@;R;48B.1NdB/Q2<+GXSMX:^V5K5fR7A+7U)/Bfc?I?F:\6]EC[FTX[
C?=)#(5:HbgYALY?X4>BQN0=Z4,ge/#=T3fKeWCJK#K()_Ue=NaeaNF=DV#8]?3=
S/S#S7d-:0#V&M+3(QD,#eEaY\DT/ea.C]5F)]<M:[6&-=gD5^BSSS)B(47FZZ)<
[YC/27]cdPg&G,@<)W_;0T,.bL[;(DG[JJG;=[f0&1\T59Ca7f-](/W/OgF#GQ>f
.[UdO3dLI]V7bQK4W5YT9W]1&=Z_-Y@A=8<N,C9I/e8T?Q)cU8W#VA/(D=DY(,U/
BM4Zc-PHI=NRA@c;ULR:6;.7,MXBKV<N4):PYa9a8G@)VT&6?7@W]?@1IL)Dg7K]
a_BaM&E2eN@^\^7IV^NV8dC6F^UbN>?/N3O:J-fbS>Df[(,2P.4cJdVH&8d]+8?J
H8(MFLa[,2N^O+:KMa2?8]G_;LJYB1KS_QQVf?<VO/7>C-S#4e\)4R^_YQSJGc7Y
-J,V^g8L2X=8F)19Y]J?,1AE+KgTEBS9^12GR;S@:G81D]B4Y2F6\JP0]AGaD=Qb
:CY7L\[CA:BN)>g^Zd9FEKM&VV^0Eb59.H:Mc:OE<.SFZ/\B:I6EP(2(R.RHOV.#
ZO-_[-)<5R1T3Q&@B3.Z]a?W2\T2\&BO?T,XgdZO61:+LST<:#^:ZJHg\I4=_=1^
XFgMH(.CFR^SSL8;/>^IEKG@[dL7ZT^)P5_f??&-JE[gHSZ86eMC&N-FdGD:)(<C
<bS,P#J7O8WeY2Oa-T3X7bWM<^g5@)56>=E@R;5(e=PS41-MP<OOS@BHgH2(g[)O
0\7:c41FFAV([+fGg:MY+W,GH5=RYJY:P[6W&f=<-<A;D7LZHKU29/WD;@=RG<aN
HFM3;==9<cO+NP>R<Sg=PJ:b;Z=\aKG>09FEAF)292EaGN+@YHQ/8,7UIX;<QIFQ
1]6gQ&=^&JD.TXZ^?;TLCdW\7bI-3/STaR@3.]XgQ^e+M30A64CAA]/\a(@SC3FH
E:4CBg7fAS:Z(JGg#+P(AVDW4?:=[(Gb(OO;W2Z9XFP,^M>;Fb/@B@R7^@O6T72c
(_DT@F0N(BSJ6@MNYRZBJAIGX\YPG.D\;c>fI+F:=61Tb>3YUF0dT5]E?I),1=aO
deJV2b7b=DX?^R@B/5a&#EPQ4@Y2H3^,.[Ug.AJ(:@G]VC<=UAJ<]:2YW0Za@I=f
R^4Pf56;T(ge>ZcfR6I+#Z>de7E2R]g,N37H<dO@J(30BPdHO\+^G?Df5/F</DB^
(PFKNQR9#^F^0[Q/\GcM2[@F7#EA4T&9(8cf8K70S,73D#^#D?/1P>MCI<@Sg(O:
KfHbV@<MNfM],EO454G,L--B?DLd1J97L[OMb,YdZGg]4BU?JgM1K>QfI7YcF2)e
HF#R4dY#^?DO];1PXZf@4:gg5c4&H:,HZMNMgA=+dc98A9fLEWR\A&4gG(1;.8DU
?-2U]@RETV/3=D32YFTV<e53bERB#P:aYTBW+GcP4GLP^H^W_7W?YM^7]J+NUM9U
f,Y#.RCc_fG^:#ccVTQg@B;9gO4YGBD\aeER.#3FS\L4@Z9bS2a):?R,LFabCAR6
K6YXU#E2<UO8#20,GUDPVc#ZWaP?Z;M<+KIdJ/>#fK]\C059PG](:aOGa#CDA10Q
dX3a8:g\>?#@<?]/7&HcC6P_=gPgQ#WcaN]36aUeIX&.G.d^7,,GZ.#[f/;aaW,c
cZA->KFNF[UWWMe&^YMgXHd#MM2AZfED##E#&>De?R37+3G8dM21^I0#:JSDT121
5-7:8NOg>9E;g4)KG8+AY-2(Q\D2/\-<g)1_P[(&2/0DJgTI7^975b0+;YX59;RL
RdVH2)GK=RFSW)N/9J-KKURgP:2K9RG8VBQ9^(6L#@/)REQb0I]aAf:L65cWSA/#
?IW(a1\;^]1AY[V,(IQ:LY/I4F2@>&21H]NO+3V[0PXS>0F\++H<AU-f6c)O<bZT
-?,3H8CTe(C4P+^BD\4edBbJ01U,XO(+fBW8\+W?b/,R_+/LLc]3U2^-^H2cMQOK
<CCbFS(]WW]&B&8d[8?IT^<@X@bGQE:@POJ8M>\UCW\_#g1)HMMPa3CTd<dP8Z^W
+Y)fKQgSe+GN6g<+>ILIET:B>34XNKcVHY\U-]]P_RDaM0BZ[K2Ab(d.U6-3PK,G
U\V-UPb:05++J+-e0)+@S:V5GVH8DDLb5OgM-5W33aQU;=_;+3(]H#7A&OOf.6E.
V.S;.Q.@PV0f[I&+Mc]cT[Yec@G,CbFV>BAOFOL]\Pf9O@>W>NOUN7J\JIG@c>L&
PK4JT3/2f\=WgBYS\fL_4R5I<K>&M(8F.>[c,FXZ\1GgaK_[FeYFRCKDeAO\MSAJ
S:,K=(Vdg#gOLg1NFSF.;F-I(+;Vb2D7FLI.,A-RTb=V.U(AZG]EMbNH_TYT[(Ng
R1]?^R9[]2-BQ:cYMb)X,^TT^\1TS\YZPT0>>6aIfYSQ(H6Ze]];00EEU<^?W)-Q
]dbM-O2/Pfa&U,>VC,0@+N\1(2FQB12F55Z>7AHDCFbOe4WN[;U2.C:2_(K?]1RA
\b;SPR-[98MTAA#La]_M=OD]F5&/H>>VVg/QKY,>CQT77\f\F:5)UNOQcCTS[TS0
Y,-OPgQCK9HJXTEf^VgTfHZgA63:4dGC8QRd(74gK7?F]dH7.M5TK.d4(I<,QF_J
JUG7RbMVLD)9EV:;&R;B)X#7D4_5=^/LA)^<M+RZ<-5JSN(#f_,gc+A;=G/-L71^
;B^Jg9LgU5HL[/YfO05I0S_B:[;[D9eHUT8O]??+CCQ294SWEMVcI)>N4bUGg5cV
C&E\cFT2_cWC^aYC\-(fJgbY+VVC+b<F\P3g)Z6;=B8\+F\HK-[OPgK1BS?=&g/U
Z11R\Q0XJdKc\&R@WcM3ZfQD8Ie_TB;bb:Ya4Z[_Ee11cUAW4[aBG>U,IM7NfV?2
SD\WXdB:)MI/EJa,5,g\&a94FA]NK6(<LC13M&U(AeJ0W]dE:#^&05A=DH[gb^Rb
FRePPWc:c;X1SA9.33#/TY]\V(8WYF+:2a-V)1.I5>F=(Oe3L;Xc;)e4\G9NTXV_
@EB#-EfbSEU/:[G:eTa92P28^a6(_&12VEE/#X)BL=:bJMW9,0Y>cZ6B-Y(gF(I]
+G&_Q,)A<&W::8]Y_V\_eCO3(g@RV/BZOG(X>=@<]3?(7#gY1-dEE=:dSdc5[.d;
C?107Zf=>d)8I+\<HLFJL86U<7\gD&JPaE;4P&+F-f4X=4&44XTX;0a2dH]T[,HS
M-0d,NK7ZUZWO-dM(F7KbODC>f5D>+(e:#L8Q25g^(8U\HV)6JE@H&=3d2)43]64
94YM#Tddg9)HFK:4gYQ-FW-\<1P;9eY23^5/fg/=2QS6a?&@I[Z\+cX[MRe(/MIa
bg@AQZ)G]_G,;Q22:5UJZ??/VAUGL1ccOH&AFg:Q34?..FBY_c6.R0Y^O7]XZD,9
QJ#2UdL)T/#OBHQOe#[APNg-)CC(9YFXM4+-W8U>2\NGIR6.9RL)?#5:PV0/fCC(
P[G>Wb&GFEOW>e9O=G#2OcY\PRM_IY>R9f0/&B.(8L3I#PON5-[R[VCUM7=JA&/E
+O<H\K+4d8AgNT]GZ,>6Y^EJdUfJVFU<J-a_dgG+_4c@R0e,]Z^L0PG[WMG->;_]
#[+.g49&--7=Q_f\[<UR[7G)OD(?I7,?AcA[dd+T^@ag3&G=.E7/(T@@@E#;HRLX
dd]0#cade\fP:IfHYK&T0;e5C<?AF[XcO@eD2<WIZL,Q00,)(f0a@\-(GA>fVW-;
a9>(F._#^[X94a38NX^#=dP3>We5-O_fZAOPR=\&f07(:^Af),,eI8C[&+MbEV]H
96-CD?[a[f.F[e?1MYFQG0,?^IQ,EG@<)OFa<?M@F/LZBdV;DUR^Ccf#US3gc1:H
RFH(]DPdMD.9f-_UFGIWeQ=Q,beTH8WIa82I5>?M;OIUXU30IgEdPUR@<5fc)c,>
K+PR/bMA\E<-[JQ81BbD2;^0.TNCJ3E07[_[]F3JP22X3+&X=];Sf9c54T>)He[a
,.-0\8U6QK(OJ))9A0D=,Y/#]^P1S]/&H<9?=[3/ZcEaD\\RaCfb7/T#CFVD6-BE
IP2WEc7Y1^,<-S1S([=JHI8S^d))EQfA:3X\d^6MLd+F-Z3_:NNH2b.W,bK>>GbN
WYOcFL6@B]8SH0@fe[2]9XT_RW\Q6>dVSCX.H)PMSWVXPH4BcH;=\KCL&b.C(=0G
D=eLDMDMS-ae[^2FZKK7[R0XSbRLLCB6TUVgbLd>J_R0)1X,MfJfRR0&TIN1&=8B
F7;EHJOCHeZO9(X+AQcRGO1dG0S]Tc+bDJBM60aI?Y#5:SZb_^)NY:,DD2BXBJ1#
.(]a7>]D@Q,#4.9&^1G/TYAHZE/O,Z<XUV)gG-2HCI>OG]P-VD1+?RF13A&&>2d9
UO]A]A_E#<Ve=KWbH3b\ZJ&Yf4_04GTd(]V[Z\F,_R/d39:TKB.WAP7_VN1<\#TN
I@VUVK,A6=]fFKMIeN2LJW[UR?=7,C7G@ELAL.?^KTHdPM,,WHBeM=+TOF&#?1:4
4^2+U/IC1OX\5c84=SUC)JJ5<BAA5&EC=N@cZ]=,Y,P,8ABLLfcGeY^JQ-CDf)=V
5IMf;gTU]fcA#FJg3+.LaD[F/]DB-UBGKQ-WIX;\&^fcC(+:,A41WY5+T<bWQ@,Z
@J24T&#/J,NKV.a22NB\_@U\>a3;K-d[,WX_&4/0U<&]0fKH0;7DG12UWT+,)A_4
ULR,C:b8NDHY-@UQf:=a&@7/WFIDW;A6g3OSTMGfUVLD6P,LKcgPR@?aDRD_fa/K
4]<A5&A5VBe4G0E4E\cO3QJL]-/_]1A2Q3g4JZRK:Z@J;&K^S?Gg^B1RMC]F1#3@
d..d35DNNYJZVXM8_P.K01?d/W?ZVNGDW_6^@@4.IV/##ZTfI0()YZG]VV:;eE#&
1RE;A^7^#F):fW<II6Q+T/<#MG/;?)OPAY1eFaW:)5,g0FT)YNRWGV3EHL<R[=NO
2(B@09G\=@=f_<Cf<I;e6+7,BGLW+EQ?)fYL)H[P\aa>L02UKBHaEGGb3B9:O/KR
M5CG8V+RN</e><c\YHFZeWM&BV.X<aUX2[UfTZ[P7a873:^EML3BKSKI9>S6E7@6
W=_bVO)ff.P#[R<1F],1#SXAeO+J@9FVbR=GLYUY^S51?EHE#LQ=LA1cL>YeV:5U
CH7+G0RIb^MNeXN)5fNZB5TG3(Z.14B9N_^7L=O@SV[DD0.CW[2[E?:)T0aXA&R.
g#:7e^R8+-6I,4H>c1CM;)TUSSA2W];6>Uac0)Gc@LfP.NA96.?POY<@>f3K5(K.
LH\_JX-c.?K48D]J@#Z6#HWUIecd[0[G,DBJ3S/0]X4LeVGW=[(C[HdZ3@=NR4IG
SJO-R@Tg:De50N64YNO_.UL:T#+A+>9.0/)-\EI3.SE]QXJK/f1-)=&Z];2Z:b8=
.^]>;;/[\\XA/eR802E)J1?5Jb&K3gI_4C5?^REAcPKC(#5JRF,M>?Vc]2_L))UP
6-Q1P)4+Z+PbU+[:V7JOcUaWb_f[L6PLCBMVBGB8PeIea;-eJYSRNO4T^46b+=G#
eE=VKX@/[QJec;c4g@\Uc)K5G0,cV:cQb?Df3g@QS#7F4Ygf>W.b[MFb@A&5(F:+
4\89=aLDWM],H1Y2cI;DVN#]aE@[e7aN&2D.f,C.cJC285;DX;,fCK-\[aB9e)/9
(b5ZZ.>CGg895AF,N)H&DLOO@6M;C4d]ZW-Y2[4G&\HV[1]]3dDL8-H+;>?K7cWa
3:FgP]A=]P<3@\)cT,fUF65O:>@-TA_Zc&e@3_Y>.UQaK,3:.M_BLLXH/A6;:9+S
NY_B914GT&[4[&\ES\3Z22)c+CdR+[<=N[9<f-[X]d>E.Yf6SgY66=A5a/G]g0:>
UN?J2P<g6cHgXO/4f;#=[4VI#+P>#Hcd]P/ND//DL^PG0d&2;C+P>I<K:&[<S@/S
(DcPJ]Y@]da7=I/X>.\[d\F+MeT0B?((HaR<(K=G-S7#ZcERaa6gF^F5P,RaU-eT
.8gX\Q84BXJ7/aEaf>[\#F\bI5[VaAYZPCFOW#/(aeO(O>MV>QBYe\5@<;@@>(9e
N?Ya[gUBTHT/b#^d=8:J4Sd2TKe([XEAC@MbY(UB[&QJFEMY0>9XULZXXWUR2CH/
.E&AGW1PNRVgT)^O<DN8OR3HR_4[X^aeTfX[Z4\T0P[c7B)^8^@B2f_P-5e?8_US
CW,e&W;\^(0V:7bTFeS\eQZYD0DW=c6>Lab):@EKKVH1We9b#g?6<XM7_)<T_cQ@
Ea9@#^_DTN>f&\W][ZLf.\_Pd<<ccJ3]FVc<SL.F5]I3:\-S<EfEG\c-.YHED3Y4
gBU;D0bVXTI:&BF6ML23fJW(3[87d>?:-SHBN+aNN,dT.I:82</47W9=.GaMPc^#
KW&H6G=CDU&IZ3c]J=U<a_bV3=H@M@0X#cBM>?TR^g[@>WaHG/I@cO>M99a496A&
a9<)Zf/;CKSZD>7<A0FdUf:TG/.O>UN=[/Da-S.M)+M9fY9dE6E2/bGdGM5P-,8,
b@+[f<N(=1^_4HYCXC)/Z?gI]bDaK4G4T(AS9MKg>c\6^HX1D^aWUBb4LAH\>/5E
eP[LME?0H@GgMNA(U7W_fc[/7PHX&Z2N)Y]OA(G#>^TP-/TefBCN[7RXW9^4-5bM
dQX&9&+BGEF4:#f,(MK=\WT#WYL)#ZVOK#c>&KdG^:C?^#[_,V[Q]LM_E2-KE?b4
La/IYcN,YMQYO^5/_Lcg4:2Ecc:2cPZVQ\e.AdL^;IF4b(.OggP[1D&a#g(0VTS@
?aFP+E8N)8bF832.H>&(cGR1X[Q\4>7;=JNK)d],LdP.;+#XALUa_+WA>G_M=]U>
K<PK&E=)/O/#&?43QY+.(Qg0;_(5=4Se=cI.DLE:Y:XF#Cb0(/N.;GH#/CFTZV(<
JAYcX5XLQeMBJ<:Q(cJUTV?K16LZ(]d)M(DI(K,<@MB_TD.,&6)FMGVW/@B#=HGM
F()<@@6OO8IMBF?LR;9#OL;\F+CK^#@1ddX7X0C[a(0ZWg&g5B?&G/GFMFBC^@XZ
3C-O@N/X6QLHUZ5S76(@CbS3J6/>94X7W[X-J[cZQQYKaD><>[(3a7GY9FRH::7F
.47ULP[:Q?+2@NV>A<AK>@<<8SeBRV=HE#Bb9Sa+QXMTQF[G@NT=L0@_9B^+D]Q]
>:UgAF)3X(Q)1[/9NgT,V6^V62:e.>@TPINE7-D01HFaAX0-c;XS@gT=T##0DM_3
MKG+4b:de3RcF]>?&2RJ<F:(99eQ,7;N4DZAI:YS/\eG]X<5D\1<fVU<5<4X]30A
.b8Qe_RA5BC7C0O]1S21,ad+S-Y5QO+T1(=I^H<gUASUb\V7=+&/CX&BD3F5TRVA
JCgLfT@949&YHO;U)QZWNBK@FI2W62dO#9;>O#8bPT2+c(g@#Y-M)8a>_,T3#^8b
JDM=,;@IIKLHBfXK:\SK19HRY13ZaN;4#1/eedCA1-@==_C^I-3PLTHF/U)\Y#Lf
T^LEDfMD_46W27#0;2T98b4IKVAT=bHb>Q7ERV<HddKPK?,T5G5DFa]BK?IXd4gF
^YP5YQJU/4KaV6ZfI078413S7VD)e512c?>1)62B(d7e9_8<0d>6Q<f_g:QPKAbY
K=K0=OC[?_L+PfV7(a-b&Y4QW+GV+JM=d_R4&,?-H.dBbW_>&e&6LX;f;YT:NOV]
0WC=7U=aT?[NMV.N#1&B_UVXEDCR43Ma>aa?ZBeg3eR:E,ggK+SDZ\.g[8eR(.]f
gN@&.L2+YLd:5<I+U:c6e/K-O\PJ-?CJaL^aSeZa,3MO?+WDG_X7@+e-QJCX;UU&
FO2)HRf;YP=MM8B5/+;XULdMXTR[eS#A7(@T##URaDPFGBU@.IX[&&04-P5YVfAG
SP9^A3<CY-a0c#/8XQ]0?U\HSbF[_Z,MTZ^]_&)f57QDZB\QL#L05R]]8c)IU/?9
A#=gRBXFQVB.14&ee,S?c\g#9]8-)8]@UDb_Z4+U@S-DD)<Q0T)45H,J]-=I45+-
?E(b=TL@cN3WbTZ&VIeD\UX^gAIg1(E7e/<LaQA=G/=[:>&;ea3[-LYU;<D;/SY,
BT5.]WF2aQ4a@)8E/UMDNOCMIZ5A6[6AO_/DVW;+IYd6CF#7>a3-Jd)CFL9#3fc/
W>NM4N?,&JP6#LYb].-.6?2caV7T<8_+_9+097:fdN_+NJJbGEII@8HZ05SKF_fD
J&8=c+QeN/8D[5/FD<S9[RL@]/W/MUN?2M(@U+Z.>S>]284Hd2;E#dED[BA6TMbW
H_>b@-gH^MV72b2E6DBU+2fA4,f5+/26HI7RY,aPMYPY@<SQ:L^C02B?M\IBP-1&
ECZB<0&If]1LQ<Bb&RBX(S_/K;?I0INWN=dR]K10#N]D6dTA/bd\FZ[V=5.\55F7
Me#:;P54=JIAN>[?&#?Y=B56)BU2T=>=<+P8#-0FQS++T_M\fB,+CYc;FHVHV52]
V1_73^)&=EA]1T#WbL6M/eZ>bUbEg0g:;]4A(dEEA[;4R6\@8S@g)#bD.<=/TF\#
13TD@)CGf\dB@XD[I4N8-L=8-FW\_>1U[7C+V;QNN4#A&gIEXB#VU>V:BU_.D.FY
I:JYb@;+16>),DQC:=ZLVNE&8/93^.1f&5]+,@LA=gH.QA73Ne/\Q&CcTVPC:SaQ
gR5PZ&4CTVFVJbJ<.3UcC+-#1XSbCWX0Qa.Q&]We\AA7D6a-]\L3(.<NWA<K+W,L
M[.][UaM<3EG_@L0cUC+-07#IGbI4UDB4b+?EAQA]\D132#<e3eH_,JW)d,f?Oab
EF3+<NARg6U2(SI0>I;[\I\Cge7Pa[]GBXTV3J8:7ABdL]e09:4T(L_4:B45/HE&
c),8X60O:-0[SS,ZV4]LgcKg\7Ab&_7XV(dUBP\Ad]FWGN3g--/_9L[2R,,R8b6H
1b6;J?^_;(E0)U;D,2Q;+(fM5LXQ,_YQ\V;6+M?UO:_R1.P67=(J4ZgT2M=b;7>]
.@;?1:#;M,FafV+[\3EY]:89\5O&QW?8@N/R\4HORY?Y=J(E/&(cZOWc,^N/]I^F
05fbZN9)RO5X7S3RH4H6[15bKS@<X;JJZ8<K:UBZ.^(TgCYOUY(MfS2=cX@CE5>&
-(aDAD.H2f;LCTQ^VP-N,D;51>O_a9/IM;b24JVd[-?61ICI^?=-O3ZI<AaYZZ;C
W/NUX]:(6>c\([2f=D:4FQ70LXPb-LbbV<+6NOWR0AWdefDBfbO&d-&Xc0#BB4eN
+;58L_:Ze)STDW:5.a\RLX8IHS>;THAg8O.3Z2>M:_KeLBG+AI&IEOP(F]((2.&M
0=7UDVgEK9T(]4J/Sc0&aBS1(ObC268EeKX;KQQbD9D7]7JH)\LC7:gO0#JPOcX9
K0T8ba7fRN(AA>U,<OA,g(V-.EK:W28]62Y4;,E6_8)<g5/T-5Q8>R,&KLHeU\d<
FK58,bXH-KNA_S5^KSN.?LdDU+.C2/WXP\._Gg;dCD:(@T:)CA-,ZU3(LKO(BB&A
SO(^+bbW6.=PeEb3IYKN#7XP92FKd\e0SJ9Z4?K-U^H?Y0e#:.(EcLS@V1d/W;UJ
R?,C;2[gDZ_B3O])+?]>dIJJEJVFT(Cg_?<=5Va.OV(3MeW;#EH)\>d8-ZFDf,4I
\O(Xg-8<MOK;;609IA^a3F0I\c1KS^()0X(17(DSC@7@<CbED2#PY17,_I^[)54?
&0M5aOX_R9?7)(C?[R)9UgF-;@JeW]-gaF?7<4dS9cB5U<P_=JPL2]OY7T^A^K8S
aXMA]V=bT)H8Q2OC:5<c6/a5FLdSg6@=3=WJ+2NG^<_OSJ#]cOD3aSK]F9bd&L4A
\,COMQ[0B1G,7SODP-c7:4<H4WZFHO6=HA&.K]+5WR+PH9dTDSZc)KR>;a&Y>)9;
OZ=&>M^,1OA80-M=G:59O,7V+=>2?</W^dca6A7G#RUSc/XR/P2W\\7Q9L6TOL;-
FL2Xf=T?ceZBc==L;5LK33?/b9S^GZZG.Q25cgT^PO:^B><PMK]#E8VVA/Y9@D4c
=X_RMKfL?=[31aa\Lc)dKLM/I_P94NaYC[D_>&1=P[ME8\YH/XJ>_#);=>=-6NcY
e8^Z8X@-<R#@8^(2+1AFY2GZ\DY-)@882,=Y0=2ZI-X[Bf<>QGfg2+8R5R42NBD(
#gJS56<RJbVL.HJ3EdYRaT.VKL4?FF.Q5/D<QW?-^OZ_]M5CUP9JY+PT]KKDcGQQ
/<,T+97fCAAR3V]5HOa5>eX2gBVLMT[aEfK=M2KgAL/<>2e<WL<IaS(SZ63JeUdG
-YcEQ.&#EfAMT41E:8eP=ZND?S.;D:#^:HH#)&ZZ-?.E6=74fP+G-OW3VbKSO2cT
4WZW+QW5ZT;7<3WQO^=SfZTHcO.-^]^SPfZ6CID_>LFBOESg@X[Sf.[fA<)V-Y-,
T#^aZR=NIQCKP5d8(Q-?>_&)GA=QARD[9,3Cf(:f(.TVSW/EF4M<VVAP(a?J5V?V
&3G[[.YGML;WB@NQ(XHMbg&Nf0EK5ASTQKUegB?FZ)+[0U3S55\@KaIbf>fQ-7HG
OJ#SU^\E@NU(FL[_.26)[P3F9OQ&F9LJ8MT@CeJ@O&,:#@QWWO^K<HWd8A[U,Y_]
;<+@2AMCPBDE8LCO:.]_CYI]I\GC?bAeD<1TMOdX+S[#Q7(.L2(aI9aU(S-7T#Rg
DJIFUHW#,#7L.Y0A)\7Z0Y(8RH@,(O1CB,HB.I2\WE2b7bg&NDNSU)_B^G0+3QS/
<8+LdC]-g@X0;R_:ZMSB.cceHIE3QT&J+21:f+5>T.OUKdIa,52+_f=g&:Ec7>eN
G7Z=^NVPP^QfM8]NZJ3?UA/PgKOROcO8-<4>5FSO)A18Cg+.H2W5:21Y_NF)D8g-
/44713<#1-LO4;7M?,O2>A(?W.5B^7^&Bgd&KQ^Aa_e=/I#;@a/E1W\S6:-9[OBR
)bCPNZBf&P8BbVbMQB5C;QccK,Ld^\c[ESB\KLP=Ge;8>b_C3+.>fDNg#P,CgcMC
LL5QORT(1E3YW85.9UO1R>_FTJ_-gS4B[SWH.=cXc3d,23)J5.F?SC6&6Pf+7gEg
=Ie[&DL\A.(WTD?\/<WL?,bD4_B?aN4NQ@GW+K@5-B;XJ0c/D7U/\);IUORe0.XV
f5H&(dD3XG2?gOJg:2K)P8?G-4cK6O(4E2DI(2(^GZa-U?M#0^,:dLU^)fZXMKK_
HB_;<a3OJG0+7-)879_)(6#SQ]FM>3C;eT7W3V(RPEA/3M[E+R44Mf;H5>5g)eOY
0#7QAb@2\bACYSLDMQ0VYVL9MGK18fcbTQ&[>O>e+N98TF-?0^I;.PRbfO-NHWV1
_>2HBYTFE6(Yc^#]Ha50RE9+]^XVN0[3>IXL,&Q\.6S_7^Cd._4[F8f/FZWcQ1eM
Y+X@5[Q02d-COU596))bP&1.T-gOFA]V7#;K?>V)gS17LS<50MTa6AK;RV:6A-,2
_&@-A9_WO=2\]?Y+a0&/RYOJ4S&Ka41XT#-J5QX_^F2;A4+=BAVP/1Bg]3W?g81b
_]=U@MWVfY59_(D-=VB+/?CcYbRBfN8SOTU]][8D<_066;-:Vc^].TMS50X6b@2g
D3I)D?XNb6a_g,D>GIBGbX)H]@IX16B<b&F5FI:S<#dL,X<0/R2DKNO.ZPRAPfaG
IO\CO3.C/OLTec?07)=aWE@.Sgc;Q(0g@J1F);-d+LU\(W-2E\G.)TCJ@NUQb?=g
0A<#QV;,b[I&6TaF8UTK\TCbM9>BS8:+@+^UQbUKg)4eW<5_df995,SdbO:8_O>5
O<GZgfQKR\A5?7P-OLK<VFfbD]dZgA=dEUF_5>PXb<?Od[K\@552M6I;/JT5QU16
W8T_WP,SS,=:OYCbC(/M+W^NGQT[>#dKgL:PX3R;]X^O9NQ>RdcAB?7D4c50->/8
?FQ5FKT]ZfWY1dMF/(-1@dC<gX=8K5K,S-AG(+cA?W1N18BU.d/7A-^QB@9b--^B
@2=[B-=UcGPaR^67c/=WR:4G<EJ(SOg9-7dB^X6&@W:)3;GL\>ILTJCFZDALJ.DV
=B6\^B8a&<>c-ZX3e\9JSgE=_0.HQ;ZFS,FYG.O&NJCPQ4aYUFDM]KGgU?&2:64;
Ff?=9fC,@,dSYSLMBBJ]0+<cCNYTN4EUB3@9X5f7?]>6\A4KMCd(AWO9YR?TZ-gB
b[7[V3/b/VT)#=N/F+FTA-_MX/T+LQ(5T@0<MaF?7-M:bfLY3X7OL_+cP@I22aSG
3S(32DJV6IMK#D>>g[LK@RMXVMZ/AYYRBCM>H\YaF55J;P:@]L3#g,CE4&H[F+XJ
\+-RIK@[,VJGBQ4>7+c\7VZBT\6.-PE:6gL4/L@42H#1S2B>;8cHbOQBGRcSBC]U
5E1#/I[JEe&#U20g0P)+M64(R=MMQB(GIUVBD]#L<e5R.:T6_YJ/YceG\_5.>ea8
_1G.J0EYAM_a/V2bVUa/7S^V,/b@J/7T).[B@U@6Mbbe=5e]TOTC)QG?eRTaBB,(
L]gIf\<?:-4C46?]9)V=06#&dg^0RR9]/0,CU3/B\8Y)e7P_.UQ6YJ.bf&^+OJ-b
\-+#K>7+gCDL++6M5/1.3A00?>3\eMCWU@E=&=GXCg[=5U4G?6QQIZS#g_I(FIYS
4EQ,=DB0H_=Z7(\;RJ94A198@NCd56W;R1TJeLeSE@>QX:6P>gT]ZC9I[F#9AY)Y
+HZL@VKXU>GFQg9P2-IdATeL-6>L9FSGe/2fEXe6ID5\X7O;,[RZ:cG+^O=F41cJ
e?#e+)H;Q7e]ef-U6S8]9LC_B<4]+H3;B3_b]8I#@3CQ7a4Q5>Z=-MV&H/4RE,aX
\OPSECEA#g]QK)f/O]eC#a4)9@E1OL<aWSf3J^c84CBe3:QLf5@SN6S#)Cd:3S5J
QfJc942@&EPK@g=G9VUbD/<NM(U[_3QAE[J<)7[9C2II+,^cYL];CEcKHBA\?AH4
fSL@KNdXXNOC:.45;QGNL>++2MaA)^AXO6_agMF(7S.C1QI)JPLRFV]8UQ=dS4=E
.8#S6\/de8^_C=^NXM60F?P(J]LA;;YO[BCYeX[]E_+SfCN7/P-8d8f+#,bf9BEY
2]DPI#@:S?N_Z+-1VW)D-M&N^1X&TE;[EfHM+PX_.cMR4&gT#P:VW=RJ?[NH\#G-
[)NQ)K^F8QTV,C7_:FDa+&4H4d6;3QKgfbbb:NT;\80)20GZ]])+PRXd5.RadD#2
E:J+]+a&TI/U?WUK)S^;19ZYFMg\T^^H(Ve(JQK#U5KZ=9a+RKaG1JZgX.^CO]&]
9<F>fY^Jg+P?]ZFV/J>CaR3U#4]@T:32L<@>H66C1N@_,c?Y-YUd<LTHBIBE]_EH
XZ^UaAQW#O_LWUZ&c&P\a0FW4&Y&5b^3LM0O^<@18ZHG;K;,&4=ggW^=_^,[G)b#
14_7M(J<GO1?8DJ;B/5:dYT,IeD35f2d[F)5c]W&15E;DOT)2=D,a:QT@-LL5e7;
MG#a\gW[\Hd(N+JP[D6fN>X[IF_.1]@ZFU;BbY::MP)(CW#EL\a((31e_MXKf=HH
<CI3f>3_^8VT-<7Dc9Mdg^Z&W=VBCQ7SR&,LbJ_S^-O5D,fZ/:b@@&a2X=9b?ML4
[/(?eMI>@^DC^\W1E1?dg\AaKGFH&)<B&\>5b(+N\g?:RK_V_TB@>Df+[]2T_\]0
&D1UIJ<[G=Be&N.92D-QJQ^;.M)#XMAW_a#@5P(4CE/9?@,(EbXJ4W+X-gR<)2TR
T^2,3;?RIG&Z)G>SE>[Z#V=-Hf7ZPFCPOLV:2R\,ZaT)PSbAP5NQ]],f/]<O1THE
7IS/Ig3S@Y/1]:8f6(:&J(SH/8+O_F.CT&X))DIA/Ggac^,+ELFP0aJbD/RC#(-Z
)L;Qb9XgO0I8E0dJB0/YL>OQDZH,1VKRMf>;1Se0+KI&<+ZR-P(QK,QDGB=NZXQB
^<NR#6.WP),:9;Afb5[<NE7.OVSW&9<(G;Q:D1ICb9>(OE;HdXLTSZSLH<2TcV3:
KD5WDV_g@)H496;NP4=P857C@?K1J[Y.D&O0e)D5a-L4(C[\3=GZaS.bXDF,da1&
+F1NYa8&+ffgPWMa;cJ]S-72::BFMe(Te_\:8;G.O@NHKa]^N>P#_DXfPLGFSb.O
#;2]@DYZgCV^AN\.84:RG\?@S=IFVa?X(G_4d2TZRKR=23;OLO0@.N_;a>69AP9,
8_7CQVegb0-NK.F>T\9a^?YME.Ab+H@cYHF>)<Q\,MI]<61\_&Kb?Ocd.^-gBI;-
OE;0AA^PW#=Cg3BON,F<0^U?X613eHH(9&1)QK];<,81(FM._13SU#\72dcV.UQ:
WKFG=#VeCaMC1=Z,9?J_becG1+K,\g]+?GD0^#.#QTE[]78US7ba0-b:G/58KK5^
D1;/YK<1D2-R8V]\H.C8BBcZBf/=7NEV-9C-feJaEP76WRIZHAQS69+F\[XG?bK_
^^YG#;0PHJW:c@-Vf69/BaL.--H]6CO#7<4_]S+:@7:AN<<3MZ@HNK+Q0ZSg2_?D
O9\1e]=bcd^G9;BVTQ32e-E;ZJH45)R@UH7:&(X6++@@agT0)S&#.a4ANJ^&PH9O
1K[]=gN=BJd<6\(2c?PV5P\2TAA4>M6KS(SfPV47?<2N_ZM3L3AQU,&EbI/=^3\@
FZ7.WfJROKHUd4[#7;bW-:[7)QX^4&9CH-FeHEcCM#JIGI+?Z4B8bKT]IIT40]RV
T-6723X@WKY5:HL,WA>^PHPRN</I.JNN=bZ>2<D/]DM=>#1Lf_VRVP4GOO#N2ZR:
UU#>C,[9a5T)/H_0,JL@G\WLD\=C4B@PK[<99[2^5gQSg7V8e7O(O6RaY?]RTC)#
YO700U(3,Cf[c^53Ne8;\a5E(Yf^O=J)Y/,7]FMR/\&L0]^ALG.8RW(8^A/,:Ue#
/6P1F)YOcS4@cUVe)66g_FU47GY#E].Aa>9Cb6d<0KCQ:f/cY7ad1:Wg[O&aWAM2
_aO\dH7aGS>T-c36Jade,T4FCeX=JJ<O4cABL3V\+<a5P,D7a[0OKd>4Q:N2IdY^
S7A#EANf)W.3F#((0bY&TJb-6(7ODE8KSJVCWD>HB4,,X&bU1H0T_:VQDdHUBg2a
OQ,0A?R[ISe^^U+&X:eS(R-:_LHJdE,G)P6(Q=4A,)WIJ]5O&c9)]N]Mbd_+W0-B
Y&dZ2)9H1(Y0Jb2)G\O5EQWBaJbNd^3OBM+H8IdcC#K20)&?fQdA+JDDf:VeZS:d
:b9Fe<ZITUSMNRJOd>c+OL;UW)6gFcV.S84;5_VHC85d6D=cSB>f#:V@)g98N+a0
O?9BMN5Ef5Z6>M_X2&BTE)f:I3]f#]0HG2-4-b=0-VWc7^H&0-1>KI-dbf,)>-4G
f5J569fc@U.M+H:_V1KbMUSPNgTI+7L/DbBKaHNCELHZW(<Ifa5gH?bIe+3c27=g
?FF2&c)#XV]3&M)J];J&=8LW=Y0@R9gZ,R5@;:D2&_S+IPLIOSZZ\ZN9Y7R-O5.S
&^[YVVB_H22G\Y?/>7_RG)0JTHaR.87BKg2GTJ_dY7]H&fZMKS66.DUaB0O]KBN3
+RJ9AIJ;6X@Xc,8f&^J/RIP4c0B57DK_&aU)KY8_I_GC.N0DC[WK+,>/]5SLWDNJ
#J?HIHP&0@PE.3-aO5K/K2-(9HV=Ha?MG/+E,(>5#=#<5c9KWFe[=gDeE&SDfec+
R#OPdVgg?[.e74I+,&^gQJ>8GJPL32]R?OFeO+OZOQS,AeU./9VAbXaSg55M[6-_
=#^5TW?T/5N(dKH6g(efAU^I=+,Ac9BD>3g1DD]S-8ERN:eE+?U4MW71Xe4b..^&
_6dZEBRIB./eZeg(\G&ge_?H4-RL=2QeY2?1^^D_Y>AOWJf/-L-?a89?7a][CXZ]
9MDbbSR::#T]G,D8_HaQPOFUJPMD/_?_5^-]b..CNJ,0+OKHDUdaeObI+I#\;VIB
c-)B.X,Z^&472IFZ3R<QZ.O@9Q((f3B?+.1^^ZSc83ZGb\XF#1V^IZZIEY(eK27S
(?DU.\2=:U6<KbRd[M;6PY\dE+B&6ZIIU/.fFRg&85LG(.#IeJ73+Bc?M[d[>f-;
CII>)aDQLFY3b2FQW33MNXEK+G:<Bc-fOFM4D\Q\+.4YA)>dPX,PS8WNY3Y_V(1&
+g)U206)K28[XT2.FCbN/I6#]J4+<KL1\4cHU-Z>^=F\bOZ)D&JI65\G<,<)H?R,
Q<Z5,afGA&8Ng7RKQ>&XAe_ac6^:-XX)M&5K^WYeUWYg+??bPdQHD=4=-aAfZ<B[
ce&Ug]Wc)M_G]-Q&9.C][&c_PL-?[;W9O@,KC#_T^.2Mf@+&YLE@)3Z-=f:M6Q5[
dK(e4b5COX@#W87d]=:N7K[+J#6BRS7?MV-d:\-[JgCY&R5\_Qb;AfGXG5NM5R,\
J?K;Aa0bE)[^&BLd>9a>-(7KIP33L@J/JEZg/E871<bP9LS@8?EY\-.=B0(N)/RA
Q_@PWR&bS<;JLgYC<=^cd<4S-eZEH4+Q_?aB6=@??N<3gOdb3aO/Wb=/<a6PTdLO
c>AK<T5H5QODa/\G6.?a8OYLDMJRULXI2-S_9Z:^<;-/&BNQ40)2ACCL9,d#T1b)
6#@54SA8,R9^(g:T7H_=g#5,(^@448(K<F9Bf;\[4WVX:Eff04[[C;GYGZ57@X\-
6eWU318=P1\^I6>^PT3;@^;C6:MB(?0B^Nba/IM=-#Z1X:JGV/R5c70bB1SL@fAF
4R@:C)^P>M?5U30K@2_A-6E]0T],7dS&JS2I,dQ;T06XeB4W]gDA?1IAHV[K#e3O
NRV?[7)J3+)/(d.KV=_-2OZ\H+dX2H/dC=P>00WPML\#/M?aUXH@bdN4]7L\/QP/
E<\@,)1EaJ3G.?BD<Y(f?6=9a:a)5#8<bfURb@TB41S6D;-6_C3IENc8G>I,WV3T
3Q_=\DbG+K@&UgDe]AVTT2BPH>DY38YW)ZW6Mb0Z-=U2FY^R0R@A;Wf.2N]ELHS-
@cUWN/[S@8_=Q:C,K1NJg;de:gU.NXN;.-HCGZ7[[;KBK7Hg53>1+8#UT3)-.&14
C/e[\<a7fH+#MIZVE9-,6V-&JL_=@GHX/dB4gV61Zc5c\?_.,ZG:aX.6PDL-3=ZI
6e^O&I8Q,e)Vb0+T=8?X3gc9^_cJ\1/9)(gHK?YVPA9)0@-7S:B0G2<_HT#VII.@
5YfSgXIc133RGU?F[Ib46(;9;.NNM@_gVLU:#4gKD.(-@+\e-,9-U,&Q&+RPARBa
=TN]PM:2NO<#SN\FfP;/aQAFOGM]+.GIT9\(=Ha)R0AL#P>#E?2=P.AGFF?WR#7c
<UUKYeMA_&D0(I4@.gY(c:R?8)K8cBS(<PNOC3eRX)L?=_PTPR-#6^[C9\&D0S7D
^b+#EfD+a_Me9#8&N@BaE_#;[=2T@9Ma9GM1SbGA8SETCY50R#<X90E6=7E5g0=g
>^[+8)GS?...<E8<AS(<5DeN.1(\/04S]+;-G1.dH[)R>WZ]g7HF_^bU2<P7P,S=
^))GHZ&g=fHS=M]O0Q0GfA:QQ&9^J1R2@G=eB?Ec>fI3f(WH>KS.S:H(JbNf)T4O
aE@c-K,2YM[L9;#SJJ(H[UQ0IP5a4;e:IWNfO(:+ESP9]WB=^^f]@0>3.^@43Z>S
JCW#_,.,O5IAX?8R3RYZ&,Ja[),S+U;ZEV20+)2)FVbbU#U6GV06NgYG_BeW.06Y
YA>BI3@f8VX&<RS=c]FKR8J)V]f&2beJ73(Y&>X0QD,8+@<\0JH@2Y2O]TRU_A98
5F1=+#C4A^H<(E\:QGY#b?6a:QU8LC\RRJ@F:MV=-E&7(5CM0Q]CQ0gYE4(-[dN,
_>968;MU(>3JVDbSfR__ZQ9LW39@aDbgX@cKA)WL8M28a/Vf@V?26<<];R8b9TM=
T9Yc:,Z+HN5HH2R44:/.>MF9ZSAU\e<+;2FdTNPECLUZH26ADBNSS1D\/(g5MR/d
RPAS95NLO\,5&FRC>FG,&WLd;MQBBZ&^=K_BaZ.M,<HOXH0PfVT@cGBO&WLeGP8D
)=VAW2NIH3-7UMDFP?:_QZHRX+cX701\=^#^da-)1DZbg\)T=.W>98_Y54T>E0PB
7I&#HG],/S(<DP7K6a_1GO1NN>RcHH\JZ3I2<^g:XS+eQ^AA\.-3De34&,N6,P@0
BLgJM&?E;W&W>T8?HMQ?0aLK5CGWbA#M+Gaf&Q&W56SXC4_D23ecd-gc9H1YFBI^
;I&7OZEW9G_AF,a-d/0dY_ZL-GV8OJAV/QH/QAS41)d0e[4ZDV;]IFAGBZ?1S2Cc
,/UAd?<O8c3V8)MdF_A(?B_5cF3M,WaZ0Q[A3.6ebTY_8fPUWd[L;^K^RH?\)02b
gT(ZYf7IS7F-F)bCEGDOA1\1UL+?P+2F6a;=N&P.<OG=,2[_#GO:U)3_,62D,g;M
1f\0M]JIU.)<##Ff)Z.M#4-TX30LdA1P]546<(+\5V2POA].?dGca40/_X(2KL)?
eNeOC(]NF(JS]>6(S#U20;U)F#I[_LLG[UFU80DX6WQ;K\NTVgE#_4/>g()#W-QV
NEdOV_N=b:A;SCH53d#R.d.P3?^Q,ZQP()@CX&b=Q#@E=N;-X[A:f[UH4N)88<#\
Q078EdMY^Q3cIaR..:_#KLI7:AfX+\DeQV_M:2?Og<<a;14#JD85AMbaETfN76V&
#WR2(@^WD+cZWI,FP\<Vb@PcCL,a.Q5@<Q<D0@SUeT=F)V#4LS-O@Te5YfXJ,S/:
E-f])8P,&QW.,K?]BH=H<F+a7(:+O&:B2_2V;,F_Qg23.2-cU<4NX-_QO-X/4T]=
g7g)JcVXB-?>b+fD0cG,MEPg3S59CZP\(>UUg:3dW4;OFFeR[<>C3aP.269\:1DL
c8e^+VB:f?5#8HW8f\NV);,GI&R].=U\fN/LY#:A5I;H\OdFM^@.MTSf6dYd@-]4
L:[T=0FCA6;:_^>7O04X8R?W]S56<[F2U7gL2Td55d)N;=\S/cWHY5)==[.LM_S>
U^.O)O5]Ye>ROc^6UNf@gGN<8,G>GJOP<+IW=e@F[+RDAQdc=H;&6[;3P2+J+0WP
#GN_bgMWG36AE.&d<b4@6d/1<S1PG0]ccMX;_(V.E&^gR2#JgQc3ReCR9a[LMUW.
]dc_ZC76dKCO9UP=#a5(:e<?V2I^V4PDLY7R8DN??8X7ddZ9TID=Z)0RgTC_f#c@
#;NJ:FLS<7:,FAZCN27.E3N83/-PH7E@192b[].[]FSYLe:S8Z)B?E/BKW:2C(L1
SD:(32f^dEFe9PES3/9c1LH\=8Ra5f\P3U3U@A&](]=gU@6MfVHde6,N2K=]IF#W
\&?5B1cX\L17NIMeXVPN;^P+;Z4O0UEQ_/H6Y-M+U>:5346g[1D\K?g)U#f75;-&
.IV7VeKM&Wfc8HAU)g6JG5_Q^[0gI]Zf9.5bR7?6+CDCJa3&[16A0FBe\VU929a.
X0<62?d<Sg:>X>48_JO6(R&B1eO)FHIf13[]ffZaG4U0[OPABD]E2f#.JK-HfIS\
?E1K_]F>GK)]KQ0VB(<;O<8FR=S?J7A9:]E2d.9/ZG6f1G;D54YRU.AW\X07;g[H
#O/78E&806eOdY;BCZH9G+fXTJdOV-[]\LL6B_7)EE.2T@-+0NN=>+NE53R<ONbV
R[2RY]&HF7C.8#ZRW@26+E,Y(63PI-@2.LWFDO/_OR[>aIKRKUH8\E0&f7)+fK7+
Fg^9g)>VgKPe2KA/,cN2/#)(aF+eN0X@G#ZF9H@D]5\,,D/K&1Te(M_]GPTU5[eF
3gVZ@Q,OLcO7e_\TE:MDM6L<(0a;GAF_9=:e;7),1agOf=@.=]7&g+PKT4KFK?X&
6.A_=CBW,.N7;F/ge4A#BXb;M79K5fDc2\[S)_J-b8F)#5M^6X=GKBIGPDRUORg;
BL(XN/>L5GFTUO^(U1YH^@Y=61=JKYL6Y/0Q](:6XS[<]#HD5?S-9U24LSH&ab+\
FFfT#<^g8a&]EPP0<?M2KbNAS(RG(aK9JSRS0DcVf>;8:0=E>JZFd4Vd:f?6<#2.
I[.&2GB?dXH-3#3?4DH1R(O7(5];5Z9]K7INIg@RTgT=J-,I.BA-.#f<Hf&cfM[a
(0=+MZ2dfO6gc?4K.8gPZPWGW)[@OF^^QgR#?:UJCa7Ve[H06PU+XQO6V\dT(eLL
&EA):F+=FV2DJ74N]ZX@f\gfU+<H8gBJ,D6e1O#aNQ&#f59F(;]LWf[?KL5EMa\\
XN83NW@7HKa6)V&:?P5ZIB8=)YM5Jc4FR,5.IdFFLDUWeX;OFHJ)_UF[BIY-#(9?
4TRWK-O_O^LfMf1=OgK^ac,8,<BE_\1LgD;IYHD)^\4f)]&LWGVYUZ26:YU5;e2\
6c7@:JJAEDbOE,_9VC+g(@PS;:)\YJ_7SY3S?<&99I)L?Ee4\^DIE836,EN#IX-F
=OTaXS7W[?K_[P)dX]=Y^2(=5Tg\b0EdN665OYA4:EGP)<6KXRaTS/\d]d+cfV5e
EB89^L,=Z>M9>,5(TMJ/@H2K2cd)G&/Z[^NV37ZbdV-4K8=L1W2_0YQS95gMfUWf
&]H\F<A\OK3:EeGJFe(Kdg88>B&L:U=#HV>B=)\bYP0K2LZBGI6MQW5NPLN@5DKa
WI.#5NFdHFdgL9<XG)NDA4^G56?\^:(V)N=(6N4&TDa1)#T0S#g9#]OHVb84+[ea
bMGHBC9_8f-ZTAMf0S)AC^D[LH)U4ad;-\ge3+4:4d.C?:7+aR7X[=:K&2WQ0T97
^,^U6[,^^bg=bSAEK2cRSM@J]a6>>G^gXLf/bH.+FDL^/X-@aN)UE:,J^0]33a#R
?ID)GM<bVQ^6XdcfH1/J)aeL&f1F89HAF&3.GO)6aa>70;W]KM(0:f15)-R-WaCe
MNGF.K1d=JYc5;D2=H969#\I/217ZU^D91U-S[U7;fX1BH(:f#E-]^@Ped?AN^_N
[Lcf/fV,-ZNF33>6_UULb7g6J:N(@Q[D]NCQKg]<IOR\<WSbW0#QUaC@Z8eCTCGS
(?S^^R56]L,R2,&UC#CTPgb0Q_ea+9>=I]84;UWI2[,YXWR^0;;6K5K)2CdKYa/C
:V-=@NUTZGTBRI\.]Ta?9&)F_U3Q1/XD>>S^b0dd47dgRe0,=c-Y&cVF,7Ng^_3E
GOG+6)[a+0R53&J[ZF_K)aUG&WAD:g^.dfYXS937=RfagBO+S-V?@-5I-).]BO2X
fcRG1-6HdW#+<Qc#<TGWI=(-,&4JG)5-fcIV[I[9UT-P01@(G4FZgK8>J7VKDH<G
>e:II.@P-ac_dW4:gRVKZ4Z1Y/4.d((>+23\YFLgI52]NQ2]@H-#E_eKA]OgA\3+
(Y84G3c0\MZFK+P(Q83G5Pa+FQG4,58C]f&Oe7N>HdJ9[J@fNV+9\,VP#CD18)VM
A/a73PWJ@HL[[+9aJ^>@O;X<1#E@G1<\/[VC]-KQF,G><0NN&RXaS]K:<PJQSZ>A
e_<IfOBR9/6#W(_dAZ[@<(O5NK--:Ac8Z_31:OPLIA6a4+&MNO\DLe5^TJQ3IQ&\
&cPb:HA_>f\DI0?.cNT<#[CP2Y/>.(]0,KI]CWG63;b98&fNL7U)Kb0\19@W=-K<
DK^)\)T0SeY+7W5R28I8J^4]c#9>9O;^QeR1/:7<6:BN,2@7XF)d5KHff,3G>KF/
/YU;9@C.4J):D<FG<2?3#eZ:5X&@S,=KZ@bSK^bVN/3\T\G@RG,g1c^7bcVJeSK5
J#W\TeVRY_]VD9E:SVQKE0XdUR,\O##T1L1G9bKR><?3NX>d:L=1HgKREJ)fE)bV
fBNfZ1?2RPD,XUD+b4CG(NFRFG_F-29FfZ8\SG^Pa2RfY_bV8:C4P&[D0<N@T0a&
8]f(2#G>g3GMCE7/PWaR]PVaeNEV3?Qg\.6dM9]R0a/AH].,G.4OU+g=:f7WKPgQ
<VK]F3X_7>UZ):4ILZG[HP1bZc;)GRF@d.B0LU2H\7__VHI5I0T5fD)ARIJ)&I&\
3bNK]NXM-?>cd].HUTSZKGH6_V5HJJYM41<4D)]da3T]HLY]Ze6<GI^><#-3>[=M
\/(ERDY7&2M\6(:@Z=_=I1_[S96BBX.aRaQ<=\7;/G6IUW_<PQ=W\;3QB^;1T-1U
J3SVG2DSeSUKGPWdPF7f85V2=3\@aP@Nd53S>(:aU\[^BED/ADUdYCe_2OVG:Rf/
REBL7PC4H+bd5.+S9:<KO2E,bHfV9B&24U&4g:;VJE2FTM0+96VcU_aQU1GbT2fY
;D^C8P@3ETfR0-;5(DY6TZQXaL6Z(I/:>T?bB)VH?I<R\Ub&?<aW^C&4I)(+=(2U
\/aN8I97JJ>^3^##@bVOI\=F]BA00M=>PXCN1.7ZL1Kb0Y+EEOLYSa#-&7?L#<gR
LPQ.QE7_A_;Y(G=;W)g5&Be_4W+>,H5d[G>=7O\DC^5CeA&LU5_?#baM;1dJH.\N
f,NaO9KR]6fS82LRY++K0<4=#d10c+LS\<?2[XQ@.&2LBId7BC6KQWfN+G&0YS8;
EE\fE</YI9>)+Ee06eNQ6>HgMFaO6eS@JR=A3+Q6O@A\==U&UaI_LdKBMF5c65c_
ed2EZg=c+:GgS07,),O-+9Z-2-/&FFS-=WUSZ#6eAb.e=[U+@8U6?a48&88#eYRG
4Z)>##Q2F,,?DfHb.+_A#RXTAU7E433L:;]@6bQERQ;N-0V-(Ng1N8C^K9>J-CKF
EHLO7POGC2(,V45?PTX3&;TbeLCTDL1GfUYQYG??<\IYBT3D5D84]BG9=6123CUX
FWOUS(aQUFecI10@XH2G\XUF::gC9=[W95_>.PSd4X\g(Z\T@@cJ+^<\bGAUON4P
_)L>gc\FB#&C6=48c:OD=];]J6M\80\AK<)PC(a71(74:#Y;IV8K9H:;L6W?0f6D
[B>J;FT?B.WT4cH<BFfFPLAKY:/0OGWNSCU-T\\R+Ud6^],:e\N;NN:7CXIcb69T
8b(3N6ZJ)N_#5S1[b:1+N1b+90+(N;O<b:J9;Kf_YSSK\-(M45.<(-c5=D1[8+a>
Q8.b]O6<e_GGb_2[CI@\MI2?f50S)RFQ?G81TOM4OWY/6)0=@B0[_@QY23QQ/FM8
,IM21SG#K9_H:AOLFNdB?8NMS#Y]QCab@f/A?:4Ke>LC01aX1]eNgS9@?+Y1W+#<
A#Y,\dVSU#WaOSGAe6WDB1ffF:69eKT9]55^-1UO^XV5([9GZ+#Z_0#ZP_Q@A]_5
Tg0e]EN[(L_L=56>50E;U;V-(.BI=:74MMdHT6+A;g,:QVGAIXT2WfC<fC+PANLL
18(7G.L<Ec#\Z;3N^Q+@0Q\#:<3L\@DL>;@=,<>6U_/F408?#2/?_Z,1,1I_57>\
.cI\.)Y-[.3gC/R8AcKQ:K-BFc5@UU.@\9Ld/c9U6H=,WUWd]THA[d=F;V>X)<e]
4YZ6eUfF>9H<(F1=/^<MG2Uba(Z7;Vc.#I_\BGUG?H^A]L&DV@DBAIfZc(\3,+W8
cedLM&U\)JEO_IO^-N5H,[;8TS,KMVVON5NE+7+/7E+ILBND[N^5ZW.cF(YK71CS
AfS1Yc^GS(dQef3[V\2.(b.,S<:4.Fb>IA7A?>UXX8@9\#9c9YM(AZ-<0:&=C.W#
EbcKY[,-#S<?KOX@e4IVf/6^S2R?QQS0^E;LHbG#4gBUUe.J(ZI+0A9b^U0H?F2;
9;/2fV,0?J@6-D+dN2eZY_gE<]Y:,2<f7R738ZeFOFA0NS&>=L_R.1M#TBOI1U]#
fE@XO5D/YB/[:+NeA1AM,3F[[)gKR8JeBXWL,T?KW7M:KJKf=:Zg:17NTC8K7A+O
NJ=d:42N@\SaWa#(_eKFE+T:Y-/N93V.Ye1H)b]JTW1/I.T6&Se.:5K5R4<-Ib^U
._E\Z7a.A0g,EabK9_DK(<.gL@-/::VOHI)8BC7ZUd4#Yc6Q^&BgbH.aa36;\dA\
ea<f<-f1N[0^W319FaJe_[f]4d5JW.+[4_+W<fR?F#XZ\NGZB9.^,81g&Q(1Afa0
/HW,BMMBW<3MES:4IPO<@g[O6,F@,^dB^YW<O,d7,6A:1N5C.KSf<F[KgFMQMU3e
KC=_/&PY9JGBf#<-<^cW+.0(SV//8&5b273T6/KL=eLT.74?R^V7Ne]V\43]I3=H
8;F[I#AN2^EH-]CZ-E<Ic9H@T<QH[VPAK(5RDH-D.V[U1N>+e/TbRTY90=Od(TP4
E?3MRMKL@=U>BIE]ZdW)&gI6V?bOKY2(ec5RYTNY,YH=_2g7NS\5MUa\)B-EeR3A
<HLgIeDfb,MX@Q#DW?96N>F5_762JT31V;;+1V1.]NI8V_#,FCMZ[aRHUOZc#6d8
J<@HV/Z&(c5dOGCEV>+CY1>,3M4UXa,=2_6c0^0-6DFa;5Ue-KA\A>9O6EMZ;>VV
P9\;QJ0\,=2c[P@bU:Q_aK,9[M_=g#EHV?[>KB_:#@DRN+=I+R7L+A+.^^,JI.CU
TZCV=AcC4e1D0B9MYNeG,(H:09,S6Ef>Se.e3V6V#;73Ed7W)RZA5fa1d:7SJDcI
cYE.O<I+5T<9/ObRJ1(N/;OCSYf,NM:+H4eA+]8IG@=SJA-YE]=b9WP1,M#.U9Lb
Md8_8&V,g7Ab1VT6a&-\a5#GX4-;Sc?D:,VTE\c+Ab)8Q1E:(gdaVc6/+3GO2cSM
Ye<R^OXC+SM2:E+SW1g>&>dcbDVD<Z[YT+9g:NAEM951PK=UP20K#aKJXe7I45U4
J@9?ML9L6CA7SQ)OOO354N,,D0;_Z7C6Gc@4;EC3?72I5L#O?#.5U5<:+)D@+;S8
2fDUKV=gQ:L,3E3VZS\CK]SP^=MOUda,MbM1K]];95R<&\H[S?W(baD__VCN]=HX
Z]1=-K_KCeISD.;C^+c7Z]Xb8V&\>(ME29K&6YgM,=^[Q#b7K^(7?Eb<L<(8?RL@
CGI#QR6#b+Kb>a)H]53Q5\f[-VffWbT5PLD=1/MJ^g9?2F>FgC]UML7VUa@g/Y6)
R.SCUCY@QOB?]#A^=1G3D#S\e(NdIg.eX));N5<ZJ.B;XZeG8\Dd6M.IZ^#S2[g?
=-\;UXU=@cTEQN\/^=1VbMaf2GN=fAeHJJ6?YeS41CI&M#W8]:=]_8@Q0WQLgEU:
JVE.957,P_a#P#T9,98,Q>QZR<17_4GBGVDL/ZZMN1:225C,;MK:\?^fQ_4\b((;
DSLfWSdQ>B1RSFT3?P+b(4)^XZ\KX3KG0<^ZK096T,cVAMK&WGRK;d2S3:^ZG06b
]@>_7FNa,[S_GMO#aSX_+(:Q,cTU<Q1dFC2#2Dd/\>(PbAF,C^+]<eAO,EQ7#CdQ
/bWKLB\1^H7>>KCSGacA5I,/;MS+J?(Y((9#RAJ,IHU5_Z.A^IL??4<F6PKIKH&#
bYIJ+?EFKC@2V4F,<D9]MRCX01c#@^e-8@.FO(F#VB,((0d[6&]XRZ55T<)3E?CM
eca_CQGXU0R<S2;@dfc3IRMZ)P8\5YISA8#(38SLST2+IH.M3)=I0W&Q)/QM>gLe
Cd47a4<+9cZSN5F^PJ1(#QN\?LL_\6Jgf1;(g&-OI(H(eL)+&(ZX>.TOU]/(MV\<
.gb9\bZ.=&@b5_ZUVL[7\R,0=#M,<6&HN&8aB(;,E(LV^D-O2gdLf2EaPb(_FL59
cO[.U1)]@5KdWM=7J18=C3d].R9Nb)YT-8:A<&4Ib<_J\KZ^NG0\R[;a(+>Pb,10
]=;dJX:VMa/45aBL-fR=<EPJW0V#:WT89KR_Uf>OEF)>WK;Ad+86d,RP\82+=SGP
)Rg[O+SOS1/Zg=42gVP+5S4eAF9f[#3Z#^Q-?[f1\De7&Z<B5adcYJJ.Kf4G_MMP
Qc>\C(BSFN(\M)U?&V;FQ-U63_SZ^@8+/OM+YJ0ALCG@+.TM@3.I+)Zd_-Tf@WA\
@.)]Ce:]>R?>Gg8_\IbXT^:6RC&7#WH-7Od;ND_.J0,f:F9:4;g:=LC.ZYObNF#Y
SW\XUX?32@2a0;4a-Dd@BbZ4IFQ]g(_CW86)f:3b<Q[:cXHfH>(.J#BJ(>_MaNee
BC;V;7#YdMZY1c-.=2K&@fF\6K7(c#Ma_K58DP6H])O5.8E01?gcGZ3F<^,B-cS8
I)cM;H6.UHR=_(.cX.]+0?9R#>KRGEH1-TXDf[R8EWUTGS+#&L?XGfQ9f&X3b)W/
JVKg(2(Wa)O24G:@0/6>.[.^FU)ReVH8=PJf^+X\OF/AHWQc(EcTY.IFYX\IJgY0
+KH;:[+&&6,=[((VO;>F48A0_NSQYTC=gV&>:Q/B.TbF&BgK>,Za&[BGX\NfFB42
J,&.Bd&I?[7282Q+9?4#SMgF^A@Y2=PF-KK86(XOaR_@\/:\&U^_>TF@Pb^b>/aB
g4U+YCN+0.LK\FW1d1BdFQ6AQ\[O9@4JH&N=aF166[70/E0J5MfV1dBL,QHT]a(b
Ng6Q^37CFM-JRU=.E>f=TJbF?&<U?c[]ga^/&GUS7GbITN\TTbLBVPgaWDJOZ+Bd
HP\YT[,^]#(E_S8R3A+N;P?4g)B0Q^35gCYM@O\9-fOWUICH[?g90[e>eLDIaO7@
^7.d>N0T&\#6DO,fY01Y+FC6S+EN1Be26SdSVK[b#859\+JQN\0U;_BD3JQG6SL6
>T9TRf:YdeJ@K-K=>J]EO3.<,gNTHIWD,^0^adV(P-ZD+Q]ZEJ<3NP7FaJ9OK1V1
F^5)+[4CfHTc;P^M#4DI_8O>,9.;M7DV)D=7CC5TEa./#VY(IUKZfHTV,G_6e)Ff
Y\5(EH7-Z,W3f8;cJ,PMdC?]_1a4L6P5\85gE7^XSCHG92+Pg#CEd01.V4.,bZ[:
13SO,>#O@[OJ/W\UMD\@bg4Ja=8eJf3EeE1^TFU+&G>/QJ303EO(N55#>?f]UL1G
_PdLb^GO@0U^;.+YZF>>78/8[)[2_#W-[_=C:e5_IRY]U>GeZVUV^I=dCgLHF<);
#gRd@J_F6UFY15[T4_>2?C),3-ETOS&_fC^+79B4LR[NBME^V71GFF54_BH\^U/R
:BV/b#]GG@3?FY<^/)JG4J(PfA8:N6fB=)1/[bSX2f529RV??^Ae+<=J.Fb-;g:_
2DgNaNCU3dGXRHc1Gc,DLeP>C?c79b6=V:\QP<WGJ=GZ\\];+PWH0TBWY.GFB37<
GBK2.dD4;TGQe.e7I1Zc)BWXJ8\.df_4/H\?;M;PB=0K0T]+E;2^Pb[/@9?3>1LW
DSbHG8ZRe\R&SM2QA?/,QCJLQA_3MKLJH]8de[Y.Q)VN\O=1V#MRI5d3W5V7)VcE
C482M:g;[0+5D#L9UH<We+bc6PRZcg:CF.65[X>1;8]G\T[/.@#BE;4QRT02D?0A
I/XP)C/ODR:[/gC)\Vc41\/<5DV_?gF;2;@6;&Sc\.L<U+YJ86PO48J5M)gIN;H:
VRU2<C6E;BE(+a]BW53/@4eJd-N9ZTML;?BHJ.EAKaG=(BJO9[W,TOCH0c=?M@cc
^3)Sd;cSa-?[\W+,;6+PC@60W_>0G\^?4G6e92AEOdV6T]:5[@>@J9<HDZb_8c9A
_Oa7+ON6SW:YS_EY]f[[^e9e:Ng6L\Tf3E>2.RXaPfe6SbQH(I3YTMQD;PGZ=K(\
g;gE9g^6a1Q>RLYKD11D&7O-0._)aX/gMf8We8ZK@J9&A76S@M>CbJ>1)6^7AS7I
,dT>B,f:TP#e@-bIFAcSbRc[,RMN6G:1]I:9Q+-60+1#b@T6YI3UPJ1#AAcdVg50
HOfSFMd#H>Y2XAL7d4g<L-eOZ8[VRUTF19^H#\7I:fXdGS_.)<5J<4J>._].YYDa
c<<=fU7We]d(SG/G,#bc[R66Aa(5]SOOJB@RAYGWH(Xd5>?[59K-OaR>/NBW2U4E
YD6]bU+8K=HB[A1_3LIeG+S6U6gX-CPf:faX4<@D)C;&1I4+T<NV,&e&d4APaC4J
..SOW/\@H<gfXT+\#L6ca.OH\gKPL)-F#1.dfgfY5Cba\YF-caS@Re-O_:+&(6cP
B?/6-;779G.#51P,HTFECISXee.0[Y7eO0)X^[AU^AfU=?9789K2O[-L=NYK<KD[
\=NPQ:(R+,?DW)[?Rb?RZW1SWS54gFI?X5R2Rcad=XJ;)(Q4M2Be&B9_/^?K+LWQ
H6)#e=<7A>Q?5RE^,K(3GcL+LI--SAFC#[)?0@)S9(eedX,MUb5(eP076b#GLBYF
Q4IfXG2cV<QF&<&&@9I\4eY>3S?[TcWM&Y:aOQDB<]/[[5V=U0/RNPM?6U=CJFcL
Od<.P(gZR&M=6f=3[XcB(;6NN37W8d.-S_Pf^FKb9E\_6-ePB-#7fT^_@303(e[e
,7>FEP/#?OFV-Kc]^bA^_]^@<ZK8cB-KE46?2OH:T</50LKX>=5UNIN_MVGd,?ZV
gXXc5TXIIL&&3]K[f19A_1?dHRJCYVHDW7]>VJIT1ADLL=IWR/e^Ng>]V.)feXe@
Q^X01(I4=>6R3S@.+6+MSWFU]/TIcc4Q^26bJ;T9)5C1C9B9#F-\TP&3],UED[[O
[9=.ZF1ga,4E\RBM:YQ\;74R4.0JgNBOd9.c0V0VGAUOPdCOcC2.ddG4D;>UR3XF
7;+W8HZ:cO,D_8,f.MS@dM@I73K>>b3GKfIJAX<PUWc0^g_)3ff;=F#ZPF7f])CW
PAQ[HG^F/(K^TPaW?)5b7KP@TI6-]G9VNC#8)TWO;aCCNW:JZPaC3&6L8:dRE)9O
HMf..0FUL++MG()\NS-(LJW<ReYKWZ7?c0-;J\\;INf8;_CU,-Y=d/]X&GXf#^4]
@gRb1eK3R>HWJb85B:VM,=QAZeQ<2PBV0/F4MYK)bVT9886&aV:@>E_61dPT/8,-
_]GPbbR-dKH6?.FIc:4X2R7fXWBGKZDGf[MeYg<aFG#e9R(7D7E\CC9O:_c?UDYc
d&:87)KHDe.957CG<H1_f(W<7gQZ+.LRe^/3eL6[3J]d,fT.?IK-R_YL[YaM./OD
a+@M>[CM<be]#8bcJd0,68@85<&4:HgNae^XRA61S,Gf<f7POW9D+fP,^9]30UM-
9Z#^HJX\XAQLZXSY=RBe@HJU\R<)gW@K;&@6M@@\U+MS2WFMU@dbK:A&.d;eP/^O
+.d;2?bARC,W4?4I_ZEW3N/2e#1S_a;MER.703@WEC/-9eSN=b:BSIKM].I4;W[7
PH[ZU(H.#VQ&(b10=8.#U-e]<A7<+K3/aZCWdIEc8/O-0fPCB][_@a@=,+()cX;2
Ve#3;K=#MXM&93;IL8L#+bN0[e378S,;?S?1K9E70#a/6JP0R.d6(/;f?AJ2-cD=
WQe/2;cGE7AWI;JH#SV=^JPd@;A,NaWO>7Lc[5]CK>.1[e9(MVcgZ<2]K3L)6#8Q
GRePbO5GO=JM[gU6T_0(7WBdY>Rc3@-OKC_A_;N\7QFJ^LM3VZF4[D7XZ[I/_=>2
E^PF<S=dTHA=/_:T]U5QHZE.0&_.([9Z<)a>KWc5XY<^e,9,^:^R3EG0_?;CXI&H
BI,]F>_0J,./94^@N&2FdJF;H0NH0P(\ZAbITD\cKSHK:2S4_PWY4>aaYMXJ[gZ\
0_(V)+LOG+<OHZT^JM0##4.a)R536G18YF\^W+YYgCd@3;;\YfY:]+B)EUfP[=fX
bDMG@F;Z^RPL[BYgHLJ5TX0I92;bNB33FS\J5T3FV>d5BeB?R+AO1Jf7C-65HH[_
)<eFa5>=b/O+JU?+?.g;eHgC+JaXWJg+Q\7\gU?Td7.V\+;eNH,#+TbO>;60fW0.
,?&=D;:M#.;ITQ+K7Nd66g]P(P5D-_G#E;IVU2K&Qe+Ec<cT-Ne&-/>D.7;UUO9C
4[K5V5C\V4/W[(_5>GaMAe41Jb2?P@]S:#29>c6MCVKIAP_a.JU.58OG;E3Mf&PD
,]_&,LV=JXMAY)/G\Obg5f^;(Y9(^CC.RXdXG+f(DRP7-04cW?Sa^/RBb(;P:[DJ
=/:f09=GW(6bPO>S9983.8_VSd05:>=77\Z?aSG5?H-.aSB&YQ\).I^_,BaV7fXG
O>gGa]O4=f;X1;317=0IU5fOYAK\_.&dM+N.d4JERP7CPIf^9C=]T#_@2KT.>(AP
)&<LBUR35OL-e0WMbdAX]K?FdHN<g(c/H_/6_,IV&>e?B7e?]U]>N3:G]CAXBS\)
Z2aX.\a_Zbb]D4=8H97&LQ9\&B)f99H/4ERXXWLQ^B4EC;K63V:1(cHA?L_&I;-f
OT=X:b/,:@-ZB]YbOR^4Q/\QdO]0a(GX8INPJKX^(&KD@UK7X^V7INWdW3CPOGAg
B(\U>EBTC]8Tae?9N(C3/>J_/F@ePe]]HK1L:_PVe.=VB_;LEI5eRebTJ_JgAC/Z
SX?+8-IB\6-6X=R#<.<0W3d5,dIEY8a^DE)HU&@-7;b.H[#c2S_;A+T9E9Tg3/:/
>F(QCUD^dTM.YHT<KT8RO)MZ7[e/W=:)8fLU(LBQYEDMD6f51>eEWS[9Y2^=?RXK
.NTcV8)/c86QFP3RQQ8NU3Y)bK>8+@P?JN6-e60<aK(1:E,LYWBJWbS>^7KOYGGI
;JU^Qe3eHB,I6/Ud>:^P;F?APTJAXc_=fA;V6\FEH(R[[OLQ57_^:d/.b1(-4)2\
-OdZ3B&F_?\]5>:)HLKfg:(UEb#1FJ:ef#>4B6U/[c^5:]<S=Z)/:TCb0&H7Z@-2
0]13#d84IeSV-\4SY.d->2Y=95Z0?-A7OP/<7@>(Nc\NB(?6PQ<NNZQM:.DS7cRe
WDBFX.KW&\a@2JC]?ALH@.RA9XS?WcBW_b4X5#VX4@acX8^](F>,4feI^M[FG1^<
&>+O>GF2+cVMX9J;>gM),+9bFfFK+>)f56Yc5T&.@6)#CKKAPMWCL1.,L&)HUUC9
bF(+0RBA+NATXfTA&?g4b_O7<W^N(#H0(8?/AQ?I?WJa0-TG7VdY(59e;KDfc\J6
<EfCBaKQIaLKJNFPNdRO/-N1fe?.X_8WI1-cTD.1+W\[+6TR0g9@#bKb#K^A3MK@
b6#9VU^L^N/7H-,V<CX:#)ZZd9KdCN7OZ?aWg4^VY+.,=:#)dZIED#\>LbT7^#..
(NHKb5[<@Pd0],6JA^gUVS(2b[Y\R@bLMA+4P,Q^L6a=R2(fMVAADM#X<S6J1J[4
24[-Q2Ha5&fFNcB.@^(CNK]7GRU]I3fHO.84Z/UbIQa3,&>^V4g)9S[)fBf_H2Rd
W,8aEQ8,>[>L+:>UCZ>Y/cDZJ?;B^0O?,]1FP-092=(B]O>_g<5>Tf-&1TU(YL+0
eD-0GA[VaWdEIgR9>d<\Wf=;C#6S2Z4V#[<Ke@7@]X17U]Y_=92^F]:S:P2_8>QC
:7MKUg2gDI@fUZXP\I?0[H,>@&G#CY=Eg@P<ITcO0IB;UF^c.CT6f^OeY6P>.>][
>MA\c:a#I:+V-7LKGNfTUPa>9<AF:23e?&_2M()S)O<_F]?F28N-P^T0H53IVJN=
,6NE9I7Q/Xg94DJQLF-gJ#)G-=B#VSBQXdf01./a9(&^WM^<g6KYb-XG+-TO75&T
NC\FZ[5:PO64@[bX@YBENBKM&;ELV_(?dJ?17QdRPS__<1?c=C_AGP8KJ8E9&QH-
/=O#&I8DC/c<#C7BZ.J>.4&=+;?0/YD7P1&:fL+@+=Kfc))D2;K\N>4^EU#YcA2\
-dHX]WE/bG^W_CP9#g]0eEEDT5^T.49T,)Jb./aN>;\QAMTFc+DZ#9,@G62=2.<D
;UF>fBD^.,IHK(5\##06?<U#c@V055LFX@BU^CITYJ4#]-]/9DRGWJ_\XDF3&&OL
EJHCEXe7cN3I,XJIRU:4)E5BN]5#?#J8CFJ:++Z3>eGVH50FV^.^IGgM/#83G5)6
D>QMJ]g,4<7L7I9/fV]IZ,g<&&+WYOWNf^4MgU_R3d#Y<gTG]L8_NgK)4&=MM4>Y
>K)AdN_N9ab9;D17^-FO7gM19LMe^IQBeWYXR4a&L1,L>K4YR1b#SP5X8(.:4^3b
cQ]E;.Z,[9E\^)?Z^#66-@W=ZFA,/D^8MV.cNP7269ZDZ70AC^CYaA8A]C.&5SDQ
;PFC5ZI5E/7.G\49P0N[+N5YdX-55<g@bb^GD^0#c-^^5@(:8X&PK(d0<E_E)3\N
Z[;5WbNJIPY^HMU,c&@dFYdU_<S@ES3HEXU^\R<UQ45PZ#gcS<6]CgK8)19K7+,:
#;WQBMMU9R9BR1GdS,>5D&N06>(5/W>BNSe?fdL)C[VdDWXYK53HR,L5)EJfL7]+
YE^)K^#?5=M:9YW]eD^1g3#.XIZS-R8L@aVWa^[.?TLC[^[:VO0IW2MD[0H<d^N2
([ZQ<63IQ,3>Z_OMK=^BZLf?Y9Oe5J/:99?RE<VY3b4L^JCe?QDUf]<gE:?\\e:[
O4OP51a_@f?Z\.3(]JEU>447^I;/.8^5PC3=DV;-)VNGO;75O2[7[=dO8.\XYW[[
17I;9F;9@DB@e3g0bW.g;2)EBQY@A,I2eCYSNVZX0Z))3\33P0/FX]c58R3T?Y1V
5\>-f2WX]bN.PIFS2.&D1@-_AR5FCR_L&>SOK9.LD5G4gaJ>SE9E:/IFV@B)?Pa=
567M\8.03ZZ=;/:JSf@Q=6Z4bd7[[9P;:?:E;dCQ@XHS(3@T/?8+/-9f@/#]?Z?^
OB&TTXRR2(A?fW)Cg2;de.K-80)a]VTWgF[E?6H+.f0D0];gS2Y>MaUGGS1#\M6B
J)Gb(f;@X/-E1R^#aBOTDV:9cOL>Z(IV&57SL-BJCY4SSVG)#(S.Q_0\JFS?g<A0
UP#X8F+O;U]V@_5(F]BLB#dMVb5=aQf&#dG6RUOdWZ\f@14HW3J@&+e:FYT?VO8<
=]G.aQTg?PPX=[BRT8C:+\7Qf>SN,ANA[?U_cc[aF6LBE&KG?C7VS(O/Q,;O1^,6
dUX6_-Q[[8DM<3/d,Sa.\MS1RdVDU-L:6;)PZf17=e]XLDZ09b:1L]-=?O-UPbIY
?(I8QQ@(bEU/)XHKSPeR>CE5b3Ld\\@:5eP(M=0fC]C26DaLdD<A0:MGS>O;/D.+
dY&dSdQZO8.<YAS0+;D(93g\SFPA5N&\6K<#\Z=-@eR16-M&^VS1>.:_ND5IUV?6
6795(PcW:GN;UHa^f-3Ae_PK<)Ae+YZT]]O)#8HQ@\bPHG,]94&VZM=BN7I26JPB
6/W^^4G=MeMVUNQ>2Y-A-W\LEWbfSRDHUf:ZdT1/V>,^DH,d4E#OD.@KW/DHB/FH
LU;NYfe4,d+>J^(_)@EBTA4/=T8/YU?P8Z8e_4BDJU<V8,gJT3(IH8O6I9QY;@4M
C+RM=&-53#2U-fR-T5WdLT5]X?POCc(\b0B8U?Q[)BTT<YNJPJ(I-6LKD/0IPH+N
6Z=f&0=9JV<YK]B]+_T6.a0M-0UZVaB/YD,/c6O&RI>;^X;FBX_]PE#6,?N(/f68
J2a)=A_:Ec;;U0PP-<;K@6a=-ac-gEP[_G9)II0;+;X9O1a#7]ZH;]?;&3baJQS-
2THQgFTHUJ3Xc4QIJ;+=CFOf?3[dI<b4XJ)D=g5<[GF;dB0Fe,VUX8+VIdf4<_<7
1]=Z\E;8@,@;Ra/)_UKgK;DP@08_4K<SdIID9G^T,F:A,fQL\MZ(XIId93A;;DSP
>VQ#;96L-EfYG^F3Z>Y8>E)MF\/g9:^+^6R1fNYdYZaQ;HN)b]Ye,bE>0c+S,>9B
E+5V&8UREUH-Y+]X5//,\86>#R(gF0=]AXSYIN42R07AgHOH6A49C=caY(D5)--_
3gL?6>\FaB8JARXX^S<b(5aDK,[DFM383P8_BSS3?>^J2&84XEVCJgdQ,<OfE\DN
\4AY-Y@3a/^[WX\WD])Y?WeHZ[MfR2T6Y8NR]RSCZ^KbaIDB#OS7>/V]3Kgee.,\
dAEGg@HNH@S9Z,4fD(9/Y;XZ9WbPEF5,U9;-Z,GX78VH]HG?YcOY,Z,cZI85YQ<C
=UfC_(U@fWSKg]U6J7<)C-=Z,VcMNO>Q?d4JT<6?T0-SJd<]YJ&84(?KIUC=-gC2
Y=R4::3WK@Q8//+d6CJPTJQ5O.WaFTQC&66Pce(_E98FFXC6.N(H-[3/N&cS7P.^
5HdU-eNAe],XPXBgT\7Se70AeNZ3JT3_PJD=Z0V-f<-ZZIT>)aV5<V6Z9FPIZN)6
HF18>fSX9M>.]21@5.Qa6-(FG.WO783UM.TNdQGOMa(]H4e6<\)0:#6]_FKR_.]T
dBJ1<58/8X7T_R#@A>HUHRRF_&5E=:Zfff</>W/M\P]04aNNCf-I,S;4RULQ+@gA
@169OO0@fBQFc47/6W.PZ3CfDb=.g529AY2DJAME7ZA+3&TUFb&2+<MD#]+5R8S_
##,(87I8Re<.F>)W:K122#fKCT(:_[++9SC\KL.9G_6;RD7F97X,9N?(<f25TC2;
e[,Q3?SSb@K9fCgOG]297749J=MOYJXB#\ZPV(1]df\aYaM./c8BcCaL5]3DX)95
(#.K]B@B12>QE)QO/?,5#K0^a]P<>4fd(@7<b4QEdd-/&eP@,=/,)\M:U(QFR<(,
UA@&.b2;MF[Pb&QB]INB4F(/=^=5AK22,(S;(K>6&95GV-Q\.)Ud_Rg7#P6MPbcg
^[<HB/I(:L>\GM5Bc2X>GXM?[8#0De1W7?POXF,;]aH=4Qb^/(RFF&G4G;?,^;fe
SS9-)4](D.R\670RgN7HU0YR\ZeG4BACMZZ)VM@]29a,2QB3GY3a#TU#Cf9f?6U2
VMT7-Y=#f+<P66PP\;?(Va#g=8NMBH\C\a@YTD>e&2GA[MCC?Cc9eZMcX\K2X#Sb
a4T5aTJ[MOG26TE6^:Q78+60@U>K?2T;g8L.XL&-dACN6d&+O2fL^3HdWQA/-C@2
HM_f=QN;C_HM4V<ZQb43gF?#LR)C&b=VZ[J4S5XOQ39Yb3T56fHMZb,f9P-bKc<?
EQ^\b<@C?-88b_J<[AEgX,PQ8X=;<GPCdgS^5]eb2N,V<RQ]?bX?cT[)SGU_PC&g
C;<I7M)/Kg@^#AO@LT7(+bB&12Ja:R91Q]-+#DHS8RDS/@+JZ6+:_=9V/-WDD-SB
@g5\N<S8FcB]S1L@D0Z-1OJ.1Z]DROHdB-_L,@Cg#67X^\Ib,L\CL8(gK-MM:,D8
ecKF#^VDPJ>[:O]WH&PM&D\4Q@N?R&2;5[EMD<Af]#+>HD-25f4S,=Zd+_L:HMaW
=ANNAfL].(a#I&;(=BOZ4U40W],PfYbeK)EOa(c2PSIE(-V3_N+R>]R?Ce@.,=B&
-M-T6]#PVNd5Q0OSR>#fe)C3.EX;2@6#G2B_d:b>e/H_cMVH0:-;cX<>(+4RL@BB
4BIDVS,7_O2K>YF16J6TF-F+6eG8Vc^BZbOI3fJ1_0Oa<MK76d-G(_EAOM3F&30G
A((#>]XEUEY(IcHU0)/5W6E/90)Z1ZKMN:Q^/L>L&2E.b#;C]E<Id1]Zf?NO)aDW
QZI9c.<X/].;&^b>>^O.ccAR1<2EY9N;La5a.TA@7;V^g[c21QQ:<-APQFZb>eEO
?P777fH5KRR,3VOOND;=LJg#YNX;;DSL]91f]COgH:0VG8>/8_AGfS-T8\;fCSDE
2Z=#^+R-cA]RKJ)GNgF#b,H+^I8X67b:BK4S\<E>(W=?NP1<2a4M.,OZ>QI:CIYQ
GSX#OF_\)QdYMG[5N,EbBb+NNf,UCd]&b4YN8KaD;=_,M-T&VSC@1V_(TMZ61b#-
NgW[cd.)8c0@f;4PKK)5f&QGI[7RE(]OC++L2)C\HTeC#Va4LZ:d,JNCWAAE.-0a
E3;GRT;Ka:WNU=U9WMQ1D^&7S;NV8RZZ-YM_<_L\aCK\(1Tb+Pe>^CL/Cc#6,5X_
@KCRc/E9\?LKDa>/QCGC:::/L-J#GX1AQ<[-O<W>QP].8#c&C+?5@RT#6@D5UE0^
@1:?^XE83]&Z(Ce6<e#4cVO@[E:^=f:O(H<OGQ\/G4@\T2[/M.R(:V3N-D^_=I1+
?;HEfS?fO1@I4L45<6,SZVSU9L[63#eDEd,Jgb1/P4:[QH(KJ,50beGW#S5^^DIe
#>RYN-BDN(\O?G@95;L:aRJaEeV6a\[MLZ-FKHB/R+017c58bg=9/eg2T80>\M/6
S\-GLb[W(.N^cOS?0G[FMHX&9[4_L(?7Ub.^>Y4d.@/a]_Pe8[7f^+DV7ZE>7f.^
_6,<W,F5.2(0G&G08/Q5DG.#P\ZD1;<>d+,;Sf9MR_;UK4_^ZN57K3&?1-C68LES
/?8W?gE^a)fcDgNbYMU<Z1ZT_)SUL?=W/EG=_]MK5Z6d;7D(X460#[5;,S-=ZeQM
f-3a,X3=)c7cd6AL]Z<[d68\-:SDXPVI9fG?e:[YB#e0>,dd7Kd+-:Z,BGOH5.AN
P5)F];eH+3:6T,_Q5)3:-Jae&6LCANKQ;@.61W63<Q@9I.XOHBF&NK3T2@H9IXM;
J&S>50OYb-1\O3DM#b;Wb8A=,Cgd>#3\0-N&d6PU6DJ69TU;DA/bP^c]c\CX6P]<
=RQD:OA,?eb_(RA]5e\TFM<CQe)6PAU:LJee5>6#U5TNPg]M0R8S,U=-3;+Q)4)]
O^\f+/RA3B3W7[g?VF-aQ,XQ&D[2T?@(W;[2YXK(]<C.@]<T/eIGW<Ug<A>;7E4[
00ZV3TfI2Zf,31T_d01>7ZKH[If9a;^S-Y\;I^[+QfPL6eKA3=9)0Ma4Gd)^5W+2
W9&R-FW52d&-ddA8MO<HQIK=,U5.>Q\0F<MVP5aT(,^Tb#W\2&YU)/6YgS8@TW01
#>F<+BML.UW(/5#.E5&Q@4CPf,QS\4R#JOJK6]e0I_DWLHYgA(>eD<?&P7@A-)f)
51EKSZ\(LQ@)J;[=(WKWedQRG]/(ZZ<b4=J=gGM/H<YY3<,XO4>?8#RR8EaE?^aT
)VDFc>c(5_?+3I,@I<&1=M^N4P/ZC\PbO_WFDW>;bNR_H<LW79<FJ]#+.9WE.Z\6
WIX:]=e3SVEF9ZMJUG>Ef<H[29<U<9\5<B^)cR2B1DLOT[H?/b2f8:VNJ4C-PK[/
@S]=SdK]\b8dKYVVd++6@<0f^@CXf(WcO&O+RW&JJ@cVF\O&/L,7L:dW[C,U3H;,
M674QPQDI913,<3@W-H>WfQ\R#:G^H+QRE[>/TZU+YdH/RFO0(XEf>B1X.0F[\A\
EMMZLI\\UQ+Z@PCAIgX^P[cYZ^\)NJee/J-C4?YV]>gUMBVQ)WWM^gQc[N.FUe=S
E.O(TNZ:<a3F\4RQ7F#CXb,(\V^B0/:Ic-L=U)-M,F3>PUUBKZJ.P,f]-;ZF-ad/
-ODF,O<?M,AS77GV(??BTceZg.f0K4;U\-339EgfL<]egc2Z4(82\3ZV,YTa-G:U
C/4A(bZ(WX]4(G/X7\f3HbD82a;Ua/&ZK3J>0>?&&;D+9PP[RU7#5XHIc(0I^@)J
6eML;/U>eBL&575J>QTG9\NI]G#L/MFN8I)NA<G037K0B-?VJFSL2XI9)bD<H(]1
3,5Y]5KBK@D2dV-&#\Gc_ge.X25;;88TU#EH\9aX<3Z14b,+b&dbb+4<e5\f?Fe0
W\&B#I/aHN^:?93]27MbLO_?,)Q/NG]0&F[WT6.<a)5S4FI&]HU.311DCc13AGJ+
bK=)NO6HM38X7X4H(G=LR02EX<(3E9T@a5X6J.d5f=9#_d#A[:5/;GS2M67^_4a3
0.0HUG+6c??RGX5,[.P^a4cZNX\W-H8,^e&F1:D3<(C[3>CeO@3Mf#I_\::J3fX\
EDC<3HX>O;30dM40QJ&/@?b]QbI/Z09D#]_H4<+]L@V1N3\7;:MgGD:,CcOM6&9f
CO0FKTI_/D)d[X1O])\a?fe5g)0HXP^Y33KM;G5:3:])GU\15O1JOVH)_)P=@:?]
>W#8B38ZaDQJ&_A5XT\)P>O78G3X#K&_JDKN2YIC2\581PGe9G>#HGU,;Zg[PO@P
439[DTP>bIR1Qee=:0Y<df+;YKa<Jc10+IN+?eX)JBF)&1_91/g]Me(46ELRZ\;D
.ZAX>Bg7LW)]BcCB<TA^P)YdaF8S_<+].CMY.YJ_0cH8/Rac5^Q82/dR.G_RL/Q-
H&D9CAYJ<>_,=&+&&],A\OK7_e]U20S&YUTAPHF1_I]JXRS_fS_+(.8TM]\5,5Lb
58ZMcGIe&)F9U74FI\bOFL.0O]J_Ec<Y^9;O8L-cT6Lb\K4Y/_6,(&12#C=:,-21
Se\0WdYcRZOXgZg:[JDTUL\=RL>gDCH[K]/3DGXHeX6MU4DM?bgR0YTQf);@G0B.
>>H&R(?YIQQe[\^5::)H)GNcTL6](.-0Zd\M:^?FEIK@U3P6NeX5;7&_+ZAQ4G]W
O]3C[DKYPL+CKXRK[?&P>Y9a/Y/c&X\?U5?:?^g-5&a0:<[TgJ_/c&K;eB@R7H(L
1b)9f:BE1/39T;^T]B<cV&\=5+7>HK1].WK]M?76\;Wf7FQaUDEd/.4SB8M]\9.8
bS0+:Id&<.B51abH2DAJ23.AT?.ZV\RE-(H?4AS-)XV)IVFLa>8.MH^2_Q[/O0d(
D3+^.aZ<2e0<\NH1H-7>a)e&da^4(+O2HNgVBgM/[[PLFYA1g,TK,P2]-F=U7?73
Wb/f_T.?6EXfeXLbG-OXC69K]Ba9>?]XNIba,.dK4=Q\<aS(J?<(@E=LA)9#Z0QI
L=(eSFGEL=)\e78N,;fCCR4HTND2))I>T6F@AM^GV\IH+])D.(6fRUUVL\P@<X2Z
YUgaFM?Z9HQ&MPbZGeUE5Dg8KeBg-\g]+0gQY9?:&,dLGDd5UAeQ#IJBKG6]Ha+F
8)KQQ&M@K?bfX?1OUNM\8Hd2\Y]G^WZGEZ2,F[>@3:Q0F(DJS>I.?\Zd[Z)R(=5M
<gMU>ce1F11S]gJ=TaK-:W[J@I\:Kf=:g3&T+PIIQNIbHUMTd7=;EDd[&B[aW+BO
<\X]U0EO75B^c4f]Z9eMb#Nb/J\_[B<J\c0N47B<VWMT4?/gW\)>3,Pc7KZ9gKP4
:F(,_C0++\MCG:YG=TWT[6&4/I9;&#X8b=\F-3SB+06;27PcWM>D8BNb#E9DWd&+
H\eX5bOe;F#X-L-W7>U4Z1Y85#^1cDaE0A18e/YgeP?7.N<NX(U3dM22,1O&9/^+
eV[5>)cMb9+:\\Q-ZB&fbX)dEX?fN(0+TdBW6G85NCA(SEL3_@+UZI@F@[D^,TOE
a_HedT(6_c#K^&J[fUW:b1bUZW:RQaX_9QP8_@9)1<<TK<,-UNPe:?_TKS.9PRC@
1-,BKT+A3@VT7IB7gY@=@L\JAc;EE6HITSS-0C:1#OG[Y4#<5N?7ZF2b:K>CQa#(
3WcLIO8^^C?Z6H]3I#f41H9YL(D)dM/B@efDM^M4<a3>^F+O417M_4B@e>0OaW0)
3Rc/)9U+_dH-c9)X6-O5ZNW\WE@?<D0UB,&KO^4af4Y;G(Ib&>fMeg311fZ&3=Uf
e-,@8(PWQLf.UY44Wga5\]PLC,2_SAS++1J:8,2D3f\LOfbCe1MKV>^=1HF8QB(X
Y<UVL=1AA?KgT8dIDf/;NS#0G(MZ>JP-+Z=?J#^V2/VR9,HA(ZA+N4dBNCYI0ZgT
-&Zd3(dTQe=;<UC>bZe9_^agMYK;^Z2JQ+X+L06MVM1eKN+SNX.<PeE<O43QLPMW
b<&Y#4\F;7agKKZVN_#HcZ\S6NKAg\EVeb8+-IO[&:2I(9-@f0YAA>-W@c5_b6LN
#^F?ATJXFF_UCHR_SNK0(RS_8)a6SF7#1#4BM_ER_IWeN:4)BM6+#8-KSPb/fT+^
VVVe1O_JaQ/,51JfUB;0&V,bgDK,+/?K7>GD#\4ZBX)4Q6cTaP94L3Tf2X3<#c2d
^:8K:H-JdF.#(&A^[HEbf,N7.-EP:6dQM[/9M,_T>/EX.8OT8<.Y3c8A+X?JdZ(K
SUPe96&fBVGN1+d>S@9X6FdMDg#U1QBD7M823&<e54a:#\Ke2I0;;VFg+baV3fAd
91?NH2--?b0f-0-CJ5GeY1<B5TeY\eb4.Y&&YH21,.-Q8[3,54,1S\7[__XIEbX9
?H9X9G18G<L7Y1M0]T03XU+ZZ#DaDDIfA3YM.F]cWXCdP[YH9:6B+L-DJ@O9eKe.
@Q7:eKFU4:S+aXEgUe^#&R6/_a?=&^QY=SHb#=?;R;.R\TE@eBI:E^f+:,H?5.&L
,(QHD^a(a+I?M[MR24),LRAP\a-.4T(X](G:=dN@2(G=\.<]_e^0TN\=4MdO+dW-
O<Z)af):>ML5-_488cQc-/WA.PPN#+d6dD8@gIgd>/D;fb+3b2<J0A&BfD_K[ZOc
;MP8D6,bR43^6I2MKN/=BPA#4V9,c.]+fZC_#1+[IB^I;Z=7=^@=[81/P/@E&&K^
S\7e[ZN986E1&ScdEOG6+[VH95FZGIYE_+C+dFA(M1C<8^G5>HI6c]TTPF^R006Y
D-b:3c?T&)I=ZRF[g.UIQ2=3M-5UI_?DPb/5f8:14F/X__g+f^,8L0WXeDB9O@+6
G,M14]I&QMgbPCM^RQa4e=-_+K@HQg3O-W(Y.CJ#?P1&556LC0+@7-?2A?L3>(PB
M)H:NeX_\;3IdE()CJ[IT#A@;+Z/1SNPG2IF_NRY=IYB3#TbNX]cgNK99(KGe:Z2
YL7/,BU2H8L_c+5EH/VV47.T2IF@\db_)2Md8bX:ZM2&G_8^a\gMID2)VA19@A@Q
PT/ZSdS4\2DI>WYaa?.3:<>8&c;&A@UTD#gD+L)PO;&+0@A4RFc;VSQK,eR[94)7
3RVESZaO0e9[cWOdL:GaEd+5F::@6Ua&+Z-983Z_GUUB]4Gc7&eHZf-J[YX]deN.
2CAA3g5W)9-eWa?/7.]^(I:Jf92fGDYfc2Q8:N4URU4&_QM_CN^E8dV7bX?g,5XC
L^O:48eFMY9&@[0<L1N-:T@\KK5D=W04>B<OE;JOZASV9<V5)E^3/\X.-9>7XYIP
<[9#?\7@KHVVK?Y^c&0ggT3b<N9-4Y&7d][ARMd4G/LRRO-)PO4@\6N@2_LCNS-J
VW>b6:>9@J)=/c@T>bS#)gE>ZW\403gdTZ146Xd<&?;a83YPWQNcIL1D-Q6Nd68,
gCE7BA/(PF@.dD@]?U7LZ)BW>SK4<I5:T9>UB&2#dYM<TGeX#7Eg]OI8/,MAYSa0
6^/6CCEVDI03V?7V8)LLf+8=>P<[((89WX:1]dEW9WJ(IO]P8\YB^Od#R>4=&6(6
UNI>3HP=HaVEc-]7+Q&V6dL)fJfaA:g^cAgK[I0IT(D.+DIHEMFVOXaF+Yfa)&.f
>b;S2UY0NVe#,,KJ;<a_D]-?&J,.>?dQ,#=f[H>7>:cCD@C:IcG0.B)R&Y2FaBDR
\Y?=eQ=H7^\Z7Q9CZ5LW[c]86/I\@)U;?b;KTLYf9=cKIT=g_dXN+b7CG;DX31HD
.aK4-56d^;gdEYJ-26P]X^3^9+d_F&A6Q#BO#R<W/#8D#d<@3J[1W;P;Gb@@]^4M
7=,VSUL_-(Z>,dBFG0SZTJd2\9GQAFWVc9(d:71TcQ4BK=-:f]=>fG;IDZP?<@M7
)_J&?FM-=Z7eQ+GRZNX;+P-aaPX&aT=5fR[@=>g]<0(8R;@dB0BA\9#L#\D(^72(
UM)P2N;AW^GEXYSDE+H6/YY]I#O=I;V?)O-F\E1f)Ud>ZH/_;XJ?Dg[f@93)_?fX
+gNDYVCQ7?gY;](?>;P]YY=FNN)CF88??<FV)2I.<N-YH1#&d03D7L>02W40IV:U
:1##C/+3c7&Y6:6@cM1=R>-1+-=ZC2&NV,5D?C\(/4d#8AC_#9dc&#RC&SX_@^GM
9;:#,[2?RSN_J?R06d4eGOEXZga)Z-\dDIJ\?TP5#d+M:/+/H>:eDX]-N_.KcgQX
KO_D<J9^CLA_@HW([KGZQ@8DaXd.e=a6L.bP1A6E0S5gVU#XQ:NB8HJT^,2M;8RY
5HO&(_V]J=\17IeYf7376&G3-,Ic7T:1F;Y3KNCO&W,UMAER81&H-2Y3TKEg+b:g
EGY\f\[^T3V2c,2F[M<3\QANV_O[9]c.a^2a)U+B&d4TI1U1)#b[:MVU2[ULYF4)
fVL-MaE7_c^JR#_V&EZf[g..KTHGO]7gO)2^cDRU>2MbF+M^DCG\JI0cA3MP0U45
eS5:[DR]XTW284eFX)?I5GQX5V.+aEL8:_QD[I0FNYSE?VdeI=4gM^,V2fTXgF3[
MZd_82;YM<SI-U-Z^5DU:54=B8T<eIEefA6JNR]\B847f1c2\=?b;QH46.e=4)M\
=,Q:=Z;1B>&TR(N,R^JBTgOUL]0e]E/E15H(2]2#E7+R:SHZ/6KH444&]PC@JbZd
@AEJBMG7X7>N)VO&:bOWPc6?HbI<^3W:0JM-5)-PC;K=7/7(a?7c;1XT9WId]J@G
7AWED&T-+5YUES5>S/,dSbP/Q8IUU/M,O#;;]f^Qd25c:?c-7/,RZ94=S+8[5_T=
E=GdK^6+0B<@#]If387P2NQYA1QdaU0/MG@FF4PO^RLQ.QTIRDZTK4Ee?BXBSTIG
?Y?\cd?02,JZ]F8E0@N#0f/Ke^PVJ2QF-6H(AgMF&675RL[87afLNSJ<7[FWA2/5
+Y??SQZIT[2e]8-@g1L2eHP+>b66;7?g^<a\6S4.SJc;dKXO\<51Jg=8G)ZLKNdF
dFL+#[RM2;CB6A:f6@-:Z:J3<M)FU/YU4Z/Lc.-e111<&(D>[+TZU>CO+CB/F_=A
B7&=bOJ8#SPEIb@bOA-)TF&WYYSV.,;H2P@O]M<GYI8P3AN[Ud9MMSJ1#J,/2;TX
<OC3WOIJ]9@a<(.?,bDI4Q:4L7c_^:PP^H=]b)/9=,[[V#;199K5d&9O7=0LQO=\
7C<F9F#dZYU)=c3TLQRP?3+PTS=2]<D+82,M2@fF39ca(=A>Pe2:V,c+]+c4a-UO
]\PE+#e2V/b/#IM/.QbHV)BM2CX9e6Z]/GbcCa>8UUHbZC&5.;7W4HDS/R@-<F#M
aP,e53e.NJZ7Xf-U+.W:-@0-<)&J_/?Z,:)3,TMGU?[.8bA]:JHgHYLN4NBC;4[:
U5RU4D>NUBOM=^K.D22I/FfIdVL\//adVFb3;C_A6ef?cgRQ9[D55<c,PZcAf.40
JbO&25KX(<=PW_5+4M_,\d:Fg#,V5c2TD-fc>=6^1#b_8O9=<5LZE[FXYOZ<E?(S
1I;]@?.@&X6_?cMK0[]KY#^5VeBX)#5--?B8:KA/aKXg.?+CN5_\cL1VCRL1=J.a
WCP6<JT93HN2f>a?;/F[^2V#8Z[;ZH6@fM)e[&;B?NQ.dNRFAGI>.B?ZDJ<C4RR8
QBdJXQE=9\KbYANKN.M4a-9GDMQ5aE&3P)3Y.C=bV>B3^T-FMD.+M\,7(0@8-@3+
D\a)(_3a4e-e4&c&1[+\JeC#bK9Y02AWE&J&6GKdgECZ\ZF:GXL7R/P/]PQ&J<6/
f13#OMV/JM#-FB[FLb\=QELQ[[gXJ#_QPg<_XX1&QJ9Y>C_7/CR6TET6CN8TD?6G
-+2DJ2BRH(cE&\)@N4E7IY2fGYV8S^9g4JZbQX=N_DUgBRP5)&AT:,6RTOOTFV9W
8=?C^9Bc&Ca.EKS-KB@HEfOOO8-8OG2IMPG9)=9/6D.LV^c8<DC-=B1T+T963]Id
OW)6)J@HN<<[GWOY\0WVKNbbga[SNPF8M1ZSYHW.QBN187.>G9509(]]R;P#-^4?
&<FXRO7TK&FCfT<15I6AI:3=_R5UXHT3_\.1G8V]+P7c/F1-:B8)\K<;TNQcb?Z&
]G##^Zb)&;EK#Z9<3dX3@UTF,b<>A=8N/W=^,J.5..TLT\&O1eK4:3UcWcQT<4G]
AC#a+T-RB/P=.b=IZ]?#+IIIF4ZO45&WCD3S\5-[/C6AP-5)5gC+DW8Fe;]-UL&A
GL(][+(0:LTa^eX68;VWVcYL+=RGZ+gUCA&V>;NQOF]\RJ1#WA6T7FNCZQ<6\G),
a7]cWVfI^<#P6.M6.-?4<@[cN?PbZUY(b3V4>O5gS/F\&\WXGL.BH\_(AQF3N&Ra
@W>AMZB3W.W;.[3ZJSD2/EU5eB1Be7-PH08WZTK]GJ^GAPSPge;gX+a#@HdgL7L8
2CUaG=QRaXZTE=a59]JHKELJVP.<4HBT_Y0Z52EgbY<&STE=[#(QO(J&.+FHP1WF
J&?0KL:XWg]gAB)YQgIF(d[8O=7H^-,S(GXSP&2@2d\_aT95(;\[a&EA-64UT6ER
SIZ^A2^=[=G9cEd_b),;=U\T3<^O2EWdDS_#221fQ]:J&=Q/&AAPAW<c,cecGI-W
3F;W2GI/P-?^L5<UB5\g0BO3H)IX&(c5MH=@e+1aCO+XR7Mg(:]_=:80;8b2,(Xd
&[=1\(/0X&/F6V<O>SPB:<U[PRKH.S-:22YY>eg210c4J^@GUOfaX(Q[E,4OMG1Q
0KS.aI;;\+K7@[[[8Z?8b5L]U.ER^W/G+YD/b;5TDAP\g^d<I[-6(OWFGN^9&/5:
<V_>OOLT84(8dBGcOfC;U1S4g,B9;^E8S.8IJMUVNGPE3GRd#MA/.F+a+/WWPbY0
OGUY^#BQ+O]/FV3[fCa8FID-KfQDA3aaWBA5PQW4da(8Za.<2?Y#Q/NE]31#IN<Q
RccY[8P[_NCUK^<fP.K>J0\;^WIZIC37Z]1L#B<,7UGHLG7>:#G:2QOcd@BV(,c8
5AN(1JETe7Z3L&9TCN=3<@Ide.>5JNU9MQ=fF52C2]E\>Pb/)MV6;)>B-+F[6egB
G)K/RAV&R]b[#cfCV+I0Z@aVQZ9YTS(@W04C=64-fM>eESH)Z7-f2H<&BZCBa<NY
;J^B/=0TY)</61N-?U_M-RgB.N>54f[4LGa/)O2TbC<eA^;CRL)I1U3WR.LS7=UX
gAQ:6LB7@[Y4(0d=dN1WVX]LF.Pg0@<Y3XA_#c_@F(ARWc54ELB<M@N,;&f2,+:.
\B=Y2Z0C@#-SX_4Y8Z[dVS)@:3(/F6B9gM0d-1A.LHReSdYZ?.CQ1ZUaQ1d,N?84
XgY9S^6:#1-65(fT62a4/LI)X_/AET.;bNL=+N4^S=a#-0B#KE@#R<]K2O_N>,SI
4(-,+\;/SJOOY_Fd/8,?6-(I?+QJ^9:TeXIC6efH6KG0&-H)a_dG9,b?/Xc/DWY)
^PJ;Y@.58)cTZ))UO)_-Aff=g[P7P\7V14C,;9UCZ1UXWKCH6\REAG1]W40Q2ABg
M=(-.9NfZ)d2/1:2F4XJC-HOaZ-N1=U^=_XFXG]Sb5cO5TPUWK5CWg#O[E#:EL/N
HN)>RKMga@T,K&Bd86a\>=P^PKOdf&>GZOaPf/RU_.H8&_H;[=]Xf30.\K,ec,/8
QQfDBH.^)^(IP9@SPQ4[V:35/2T+ISc?25X\DI/[B^]@ZY-=IFa0L1Y7EeN0[;XK
I/&29>-3dI,4TGS9\dcWOc<A[:cW(F+2?))KQA.IB2,6JDE5(IJH[J5EE\a-A4^H
D>W&ecBeZ8WdPT=K#aL(6-PM1/7W[#Z>SZeS&3eS@8DcFb2?A)V/8@c=S?C4)A]P
);B/MG]?S0Z>.\ESNLE/XAd/L?^fEf[)_,]8S.C_0DP&9Zd4):4.3g]2:W4YDB[Y
(_W;G/&2[<eG.e6.AYc\KUJ[ZU?NLN,Yg5a>MS/K?<NM):0g[1I:]e_@_Z-NX-a<
dG@faN72804R6,AO,_-g.@0M?U/GBU+((K62MXV#VE>UU8d?RVWQgf<Saf0I=(TN
/>L7+fZ\bB:KVNfSX#X;FTcW;3Z[VNK)6Yg;G4D1caCff@E&.>2QU7@66A:.VfKe
<(_06(?RNLCe754SIX:J>V3eOO9820G<P@-F38Q5./#H_eVP]CK+g>LR#WeAW;&L
2-#40>Z.1UX/D2W,=Nf#K6d5Q:;3P3UT0.Z4b@RHGg/<B.f==]I.9]#I?DM(b9)I
&05ZGcN[R<.J[RK@bVB_GBf/J;bR@)#MTDKDgCAMFZPM[NXY#.I^@6XX5[4fKP0W
JCe9MWIJe(L6Ld?FWSHF(_eS_cN>M?/-dW/NJW&,c@/_:RMc1R;)Zb),fTRf.^9+
IE-7f\_49O\S65]N)GRf:4=0ge\fK]g,&agBSeY^SFf.1O9b0,&G1+D@(6EPN5V]
Q>?@M?-/;JHM/c@MT28:8fSd3]^c4/:b]4,/,eT-(CIPOA_,<,/\YVf;cM3YL2A1
g]3Kd61HfQe06gd<F(9W2?9G=_g:4FIb]7a?U_A</8CF8,g\:E#/XXZRdF3=E^O,
)4B(KGW2/T.2^PUf:0ERB-SDd)JR;-_GFg]I>.?6Z,1.&X5G<D-57F>W-^eP1MgC
9,gO-4(CPH)32#>91dF(K+FCT&(4Ca[OIWJe7geH?<Gb.8dZWS-XDR15fCNKBDA/
51J0d16&X65:<a@^7K9g@M:J9TGaK[FBg_FP,I];3^Q[.^P;EMU/9F&=UC)gAU_>
\)2)HbK-OFc)O(VV/Pac576/_bT25_@CW/-]\_6<-\F<1G[C@8@HZ2M(::YGf9)9
91KORZ-XT8S4MSdS1]#F)a^7H[^LaD.I#?CP0AYg@EPP0^GOd4>AcU;:e&D0N@YF
5USOS4I3RI-O&^CD]LN/[:Pc.P8DR):WH?>7<a#QN/106KfeIP>?<07BQA3LTMTO
F]d+6Ng^GEA\/0e[X(<1-9gdUOUMR;92@X,86?ML8#D4P?Z9fGW\(FJKFDMZ&Y+]
4O,5HYZ4F:a?Ff4&XVN(f5Zc\,E,3bQ[NH[/4CCAXZGJ8G3fV+-Z]BeBfO;AcD<(
IFbJB0)&_c[OVE&UP;)8cG=d3C?-G(-)KTYb=E)^V-/U>Hf+B;9F8H<(b<-g9A<G
Z(=.J+[B):CPBg-1J_R^ZVTN+Wa^;_N@Y&f+dG@-5PCLK@<]F-=FR)-QGOP6W3=[
:.=Re@0QDf&_L3;We2fgNDEUO7\K#S:-<+R1ME1V-XZ^M+.WR(1(<gcGA?(9V#QW
g(a?4@eZ<47_/M1=??6+5E:90_BJ&Ba0GV#J5:BYO/2B43=TJ2bH#]V]Z&V@.)^6
&a>7Z2T.?=c?P+THCN<MZY?P6Za:DN.\H515./Ed+/+PM<fCW\IQ8>,^9g4W8K?#
d4VG^@D/C=F58V]UHKE@_Y=[91HL-Q<TQI=1=7;(f#@+;a8>ODWUaUC>fWf^dSa\
M8Z,d7).#aCM?9_GU1<N[OO>dQ4gZ=dI>B4YWZJgQ7^U=I^_RLDJX83/MAIV7Q9[
,OZ+UIQ25&DeRddXf6W_J]E&\U1f:d-F(VadY;c[PEQXJS_;G+\[fB1C+2\,4+]4
GOAfcDDHX10AX&O#J]:G:M^b.]<cO:XXgNOdQ;[(@L6\VU=(6bHeORRT,0TD:]&@
,:Z1-P+)M3A&])I\=>)#0K(;7eNF@aUR6OVOIa,<V.=[=_?4#e-Tf?(AA]>gUCL#
S_c_#gTbWZ#9)(cG?NfG/\D[7b;BZ/.f;&8TZgeGD@52ZVV.KH#OHcE5[M>70N)4
#0U12=>H#g09e&6_^HGW-91R/fR1D2agR&H7d?2>b^G[\;>MeL[6HdD;SaeG3C/R
WfRg#GHX6VDc+?3\Z<;-;=b:,WQPR.0TJd_/a<gC^BcI(+Qe(-R]>3fS3ZG8V6R9
5T]5Ib93SLF>IZ-ge@IJcf\A]7#(#U@\Tg.V+UVdS2BSKZQ#/?CEX-_FM)93S0dT
OMFgJPVVbSS:ARC_@9b)G.8[&P)J1RJ].Z.Y1&2LBY@.(GTL29Z&9a0ReA+=9Q3Q
:FfZ&(EUF(eQbO16gb<1Q5<31a)?6_N0>#MGI>LINZT0K1E8HQ+Z4YO#,N&U7)[0
BLXRKGEgHP/4/O;YQfV^5<&OMY9+WFFPA2:g=?a1L:J).3@GgS;/K-7H1<L0L/U.
NT?;Z5<-#<<bH.7^XH&F@(Hf)O@N6XY3W/R,ET8M(\ZM+-H(<bVHJW,F>1K>3bf8
g8#158)W#6HVVDg.#6,6dHXe#LgY73/F2MJY_:IO#ZZfcb]R)92)&gA#7ROe:LX=
R2&UD:Y./4O:H(-#^8_M,G=SGGQ5eBP[D,/J-=8O,(-I#0W#?6S[&)+-609TW5#Q
b9ZL<b/VN@R3V#D^F[d]V\?5E01DCAHPQGaVJO8IC@FWge)4YBC\JL-L]^c#I\#_
PB,I_UY?=6Z2Eff[&KC5Bd2)I6>C35a<CC<#c0SDaRHLb7C<FbB3c7MD-gSNH7a3
<bU44]@cCK;^[4AZ1N?59BW02:fOV/;7Neb]0@./^39Y(c)YJ=c;DJ2;f7X?OD6,
16Y.AF3eCPV.<5^]5L8K7U>KMW(ZHB[d^_1Q3?_@3N_A,1-7be_Q]MROK_9b6#N-
)=4^K/af55M:HB]-55B@=&NM<&UA68e93(>g^L,>(HcQ>R9)8FR(_a1./V9T=Z\E
2@/I4_Z[N;GHX6O?-M;V>5bV^^R=4&E6.?\7Je>JLY2W8e7:/dFd&_QY\CZe:.WV
BUaH^.QefMG/cEINe1W].8+E&^d3PP&c^OAe(-R&c-C4YbWG=d-b7:Pd8M<QDM?E
;>;83LNbD.W9X,9=gYgBa((;XOS;)W-;D2]AM3JU><(fJLe8Y)8TYZ37DM&42\C8
92b)QF#EAQNMD8\L2A0/NI_EW]LRX&8)-/;CFM:-8K\JfBO90[,US[#bGG1#3E6K
fC^.;MK#:1R/?4Ld<cR;g-N9eFDA+RF;STH6/eB\=B&M)F_F3M=R44)C>&DM)9)=
b\VaLa_fZ#eZ&LO.TX4/X(bQaL@eB<F=E=71Fg?g03D<d+QWMVKJgeX;ZPc/b^.0
EPZI93B0<UJ4,b&_gUKZ)[gZ&T+,U7_(C25250,+:C^Z=<b:C<I/VI0+a3dI0I-K
IB^bgY[+G[e1RH/?4T9DNJB+<DT;AERHVFgOZbBN-[/@XRdUY<;=J?#ZE?1\;d]E
F#H9[Yf5[3c\L(YNGU;0..BWdO^&Q).V/][JS[]YMAcgCPH5aZ=M,^^Q;J+1G#>6
)fb?K8B@>:26e/5+\P<Z=-H#EB3^3:)YH1P(Y7Cg_Qe(.<HQ@&<5gFX;IV2Mf#0_
G1N#@X4W[dVI7L.ULbKO(1)T/@Q##M4Vb:.\?S9#XR8IWbM5JCb]5F#13\<&-(d-
LS;HO&<8?@G5934FQb/@SX4/_QF#.2)f9_H&S-_#^^3O3]bL3CdC@3b]fIM4VSE7
>(WAW@Q9,V#VOdIM;/X]=^8<90>&[/83beKF.?U+A-N&IAF.,bc>\fW.Ne@)gU/a
c6\,@ZAG8&^[[/P]KdAT;CTe7dZ[-d0P,#REDZ6LE9FgQO8-bL<[9(YUSXbF08KS
/S.B97PG^7G13QPe3Q_)6,ENM9Ga?-++G97F(_)g)L_5<FO9B-c=#1I),\b49;MZ
cS@T01Y06O1H.\BAK=\RV=H&WJcU::A7R]_0@gIAN&fc_S/;MggOXL;CZg@))]Da
=C1-d(E=4UNX4J7JKaE-UW43#(?6C:;^6=F:D3fa+Ma@(>;S79=8U_T.8CPJJ[N0
-YL#7XagXc=98eQfN.^gF.,N:\g3_&0YL/Q;L=/JBBQ#\XKf;7YEQ:S[f[<AZ3f7
DH-=6;UL4SJ_92X)7&a\F1CT)Y@+cNBHcMd3_H5f5XL4d^\4#DY:dPH[A-M3V1,W
=FK,2GW[d5VDKX./9_S798RQ(0U:3.;Z:dK2[LG#BS?FF@&IdGdCJ@OD4#U_#SVT
2aAA,HV>g?+e0@_)S9+)f[,=NR=^FG5ff#F_g_6&502I]?X+A;cW/8G,3:f@R5?=
L5B)+TLIYaE6Z[B#[b;f3DC[X)GP-aAXVFQYaYTd[AIU0T97.HdRPA1LP-VaRB_g
[JSf[3=G_V[;\?WFU#35S:./O/H+^&Hd2^d^K#^1^08dK:L+b--5dFBR[EbP1W66
HW\R.WC0G2b8ICD?#PV[5?_e=Wc,O2HMabc3C>J4>OZ-6<;D0FF0+5WVS2P3U,H>
1SC,T47LgOEc3?Zd2g1G;fJb/N,IX))YQ6&#\);/EH1;W#^+B=((a7#N;UAU5dYd
?IR?<-UZB41LTG&^BK59511S1f9GJ.Ed]VTV@GG7HS1L1E>[I&W2UWJGdPeZO0G4
<>PCX5.Y,QZWX8X#:1RC>609MTJAE1)[QWLK&;.RS,G3N++@_G;2.):3Hc1U:Ge>
F-7C)Z]&[aU07HNTS=Yc7bS8R8H_@g_ZENb:bH[,PZUIT(>,^CP7SbeHV<fA-a=V
>2LK#:d@&2KaJC;/>8O6DCP0cb?Wg[@;YX?UBZOO:([PG1/7X_>YI@+QG,U(V(4^
8_H#TYRKOY:+X>\_^#)6;)-]5S7;)YY.A-.U;<(3&RQN>)9F<,VT7:B2?ACN9LA+
7EPW2LNQO8J0LJ@NCK]R1Y=ND>BCVFGe/\bN9>4_:,PC3b53/_HEe.67O7f1CT4@
V=6&+MH[6b]GO3RB6=]Q]=DUc\G:J9aS^:2P2]H\&f6+TZgACLO=9[&;P]/[0]T#
VU)ACL&OdA@ST3L;GP?X7)#).g,-&IUfgF>>R+W-;WIRE96:D@cGU_.MOGgQS-^:
@d.?Da.J72E:6/[EA)cgZ5L[C9@JS#P\T:C(c@cgG5A=+fQ@M4F5a3#?\AY?W=.>
U56P0V,7RZF+A-<CeOVXFEK&5]>A:KTZMJT,)IYbMY>RPM-cH\\PG1<(]5?GG;e:
P>(S2L_:_#J_V7dXHd,g@eCX#L/X/7IZ>76QQZO^+6fa,Z(]U1-ZN9/IS;AE;0]3
XdX57K>NZ^6Ec1WU\3bg2.17,YPZR+6>A(52D_Ee_Aa(E:;b:We=:eZ/:8)P;T[5
F#EKKE;QD5T338F-@G;U^_GW]d=dX)L>KA\XOUC/g/aY-[@XI=<J8+:O/(;f7eHO
O3S+]Df+\CO_:]_.W/P.>D#=NID(B_U]U0HMV,4TBK)eW1Z]YDO66(0bcN).30-0
;M)A20OedbWBACCX_Sa)e[R)HG5CeeZ<>V2[2:^4=)>=.g=8X?8Z+#/K7&LD1;Hg
<D[Ca9QRCcFg(EHXgA;@dMaRDB^MW\AQ=)[[a=NXV6<F0Ra#WI41GDF;&TI&_&O]
>7:#U]?<KWSH8B8&P>.-9-R]1#]O^g.&(S&(+,7+KTANbebZ-UAC;bB0PbQFD6V&
07.N6<OQd9;FWF]5UPOHU70^g8SeU5DTD.NXEED7;cS9Je?J1(6_X)\8F>AG;56W
=8#_@L]W1Kc@RQJOE^0PZ,F;GYV]W3agMY/W7C#FdSI7V6[70Ig4Zf::;KOR1#8G
Y,O+6e:VMbe3(3MZg:/b;JROS8=+eB>ZH1H9V.Yc81:;BBPgW2f9.6Mb#6D#(dLH
_dL#dCUdN2SMP7b6/.(0;5]1X5?(OZ#YYSK;S50,,?2]+VUP,ZW_1C7+J,dV4fX:
D>5[4W6NXf0b5EU<G)VC--S.Ef@8U,1fE^^<-]&4)aG>aBSKB3Nd67a@US::Kg9Y
L6f9(X)G,+Oc2cfYf&9.&F_XH^M;AT#Yb#.M/RgW7N5LS5V5DCS7&IC[\,>8NF-I
BO(0+L?)eS=2JO6LZZcbB]JE<R^1e][Y.2?Pg8[/&(-3PK522OAc8YCcRCD=A/RR
cQF09OV(JU29Z2)/FKH3NVdS>TGUab>NWg/3T&1SJ2RL@40KXK=.bCAG&J.:AP/A
(;Q(6Da?-7_e:-M1;aR>X.)5J^[BE/^C^QZMYWXNWg6U,:,3]8HNC&,95Q?F\(S(
WR51QZ8;+J=7^4:IbZ&2KY-=E8:K^M6B29BK0ULX^DH)_:]WYg\<86SJ607Y6?U^
_X3C6OTcZCUK&WR^@_5e^[0AFE5dBg:O>P\:AG+=6#HY#bc(b)W+\^;cLB#fe?YZ
?gM?,U3H\I0^JEWU@_R[4ce@87d?:#dgS][Pc^_=5Qe4P_aS-N.7E5V;0SVQ^8Y[
S+bNT?-9ZOYgIgGEDPLc:cU@E)8AE\#ZU/HEYJJ9ACe\JO6QYgMZ\CM#SP\ZfSL3
7G@H-:CW)c7f_\a;^INC>8HFT,.HH5&HY-<16YB8.O58EQL_H[AQAb_/=O^Y7&IV
6,Y2.UeM^6=c]1EU\_>D?@CdQZc8aaC/?\0-K->QbN60.V94,M:4GB5bXAU[6g9P
bYJ-N##^fa0bHX^EVAV@OP+3LPJdHGNLfSFC-7T2b_HfD3eFP3I3U2-)ZX=2f\B#
B<g_cf3b;c7HXC8=70d3dV5>A#5Q1UPXRTQ94dcIHcS=J^6?9cPDAXLSPLQ6@eF/
/-]2d&?f:MTdQSDSQ_Gb.,QX@e-U&NF^e:4+JdW?L;]QLNH<&7/[99>:F>Xd9B&W
TAPV@7TH^L#4dJA#Za91M@T?@WcGaO^,X?/K1aLY4P?R\J1(?-+GFeL8R\SR^Y\0
eN<MF4B3aH]F56Cb1R,0bU2CVb<aR5>?T41W(@RMdgCC<G<e(]JIT=?\a/(J=FYR
;<\MFJ5\#_a1c0J1>XdNc#T<BWXUSdF<7+7_gO;bS#-R>39WaU?>OBQ8>#T^QC6O
KFX_XTF^G\6c(GMQ_0CaK.[7e(?beNJ4A6[Z,O;=)HeaQX5c<E\S,+]S+U5QR14U
<9QfAf>YA;Tc>XLB2=LYFMT/W8;6D=EbbdI@F1[e:DPfW#V#_]FgD[MHfSM,C.f5
2U/fA;7R53I+3f=8S5LI]B)CA6&2[U-a@5[f]Y+<Od/SMFgAJ0&)/.?_;D[>X[^R
<R#d45WfI&]g/CS:Q2eB\=JG2W+X4f&Ya#H_#<d?M=(D;ZNCR1C()]Of0AYcJXC/
Nbe\gJ,+26T\#CNeYVTd=#(TE\V^#TVH=+eBVI@36A24a9(a\#Ua;d^V8b/fI]-Q
_Z#g??e6+G-F)b??UC5DcV^Q285Y)2UD4<5F&&KVC)R&)3Z;VX/B^Z[RSFV):N\O
e=ePXT1+4C1U5:&.Mf@I(&.=1e=^&QRIUG>L9BHC3SUHR@@6<^Z1VEEFIXTD>;DE
CRSVVbC[.g3fPaAZ?2SaDJdN4A6_?W4YfGV#J@C3SJU](=YKSU?eCH.<V[Hb,JLN
V@AAa/fJZ:(\16)]7FMC)76b2=/?>dSg/_b8QS-]EOM^MS\feXH33?:]C;K8?/Cg
FH,?TS)<KMSKVebI[AJdDX\19CW@1VD2)OC314D\N&OJb(C4@F[F;NZ9DRS6ZBf7
O:KJ+ASbY[E^8.=3)99A8.W,C)5Y@21QVaLAD]&b+WCge+)R2=[9U-#ZA=:8P6<A
L8g]#6W:BaR\;N\[>YW\(#&[U?gFOT]SMM:D03ND75eY-_\5a(F1ZCW?TeY^[-RL
N8e2a5Bg64.,9C:cc\b.-A:cOBE3e7D]C+<eL?GMe[&Oab94</ac;BaYQ@/#6(W(
b(+_](I]1ER]dZSF68AO#g10a0J1H>C##fUg14WPaEd#LZDf<IZT0J5PS9D#(5d>
C.?N#-2H)9+FeK922W-;-P2##5;Y/I81++K[)gA7QT)\\Oc>=B,[&8-NA59D(XcD
[R?gCEK9OMW7R)ABU>8Y<GB,Sd-Tb19b_-9??=@fKTIY@#>=Tg]Ng,cSEJZ&W5EO
>,RD#6C30Z&7(44^>5gG0ZB>/?RC/]E/AHc0I;(1C(G\UFX_aY+B^=M]:\GeRfMX
5&I7S.TN.G+WYT,M0/^0R1c0VL:KSJD]ZVW12#7\VX)G-?08G-]7HL=&R]F][T#d
@#6H-SF,3KU)WHf#&Q//HK;OU^R^14T&3;c<TE/OR3X,TIFb_1E0fHY,>90:WGF;
3DP/#eZY-<gCgP2Vf]5gb:&/:c1_A#fC48_Bg==O4K9#2Ce]6Q:Sed=5:)_L@6AR
G:@bFZ85K),<NN@Q@QI\RRJ.J#@T-G8_]8cLA\:5<A2SG8XD:<O+/9+L2</SR9N,
Y^<X[4QCJ?C1<?=]Dd3A3dP9T0_8UX#.78)4?80#PYVGBbf(@eM2;/8\aaH/?c?:
6KK57)WKd3<e9-<_d[cQ=)1AA<O;@0#8X_+?+HY/0HMVY2,?U;a0W>(.Ia,-US,#
NFC1WQ7Xa=bfWf[\-UJ[gOYD20X_01R2?<COQL=bb1dT)&X#S&&9.56fX/XV^4JT
(fP5d9FJ1PcR/F,V6GDgD?9[f7-:]&4baUD]DE[(Xf9<(#6P@#PQ]XPb,QBa,N2H
6L)9<F8),dGF;J;-Z:47R-gR/bJGa@,gGH<gK+Tc=.>#KVAU0O1N_W7(?<-5X<5J
\MESf)A1a/R1bRS)Ya0I)1<c3d;BDL<WQC,RZ86Zb#A)+\DcS(M\ZQa[Z/,1c>:^
APgMK7XXKW+H]?7]T?Z+>A&UK8I5Z-//CUCT-DW__9\IKH6M[<L)b1Y+a^Q2RA51
LgGB<K;RLEcWg][O??c[YKX-c6-<deT___g;,d/M=/TT19MWfR.W8aEW=KO4bBg8
3T5QREVbQLN6TSQ7Y-B_f5IGVJI(f.TS,+;;3P]RDJ;:dbET8EgT&@[KVDKR/N43
2-BFKc9XOT>FHbKeWVd6SFa;>)HcEeR6acUaCG8d\^ZEIIN,K944=9\01R?6^[YY
N.B;780>OcZc1gHeV0=WT7[/]_SIgW59/eN3TUF-L;7@cDe,4e60CM;99C+::J38
#R4M#N5Z4TI6HF,@#;N7gWZLP@?0&7EYbL0eQ9N/6=SO?3HOU;+Z++4JN^EeGGYd
^N;0>36CcCaRe-GCZON=(@)+/ASg/)1fFcS&dJJWDYHL1OO5F^eI@(+,](eMHf\A
@:T[+FMfBP6DV2YZPUMSaO]5E+eO7VVJ-CVR<\XXRDB8C6dOMggCd3BUSVfZ]]O.
[g#K6,\:=N/g==E>47R0^UTDRa]3c(+W^#XCL5a^g\Fd5P&#^d5O[416T<438:RC
OBRTI@7ABfFcZOT6D+-QF5@@7C^c6#B82.)<&LY(4ZGD1SZ[EYO/Y^)fZN78ABfJ
]=3Ogec5Z?R+12[Of,aA>.DWWMEAW2^L85d-,[S.-\\YH1<MU]WA-T;cg,4&\D2F
1#MDE^P0X(HUI-C8XQc:Zf=DVaDKM0UQccX1-BZ_NUge#;,f-AU1&6GY,W-C_\aD
.WQ:\J_S2@b-N0R1[9e&<UP7b=2/X8+&DL)Y4S_C6_#9K&:K-,H=A]\=>(@J-553
/[;EG2=_Z07_YH_Ybc1^b=H,<eYVB2+_JVa(9\JD7cac0MO&L1;G7bMX04OL\7>W
GZ_5=3_ZedJMUeIJ,8)VXJa=VQ/04@a<,McU?DQ?)@K83?TfWQ,PE<XVVeX7M4K/
4B:gW/QD2fN^?T(^)]//S3DGAF9VZfG]13fST,SF:[57.OU^E8BGR+be,3C_>gL=
W9B=>gY60BG=?e3Y8:P\Dd8DUf1a_K0a3EP1GO6+N4eOB^YUJ3XP:g/\LFaFLN>F
JC6NAU^4<=R1]feE&._=2Y1^.g;>VYH:b_[BEQ;(S\A-W)b2_TIYR],L;JY1.4P&
TK-14P9];/:<WF<Q18<IZEe9@=E^g1Vg[b6f,FHV;Q]Jb\,c\)HFZRg)<,=](HQe
5,]aB0E=f[;&^M5DKM61eII>1EL/1COD,ZKRY8<1+-agd_3+OJ9&:.gZFE-7L6>C
f3M1#[>1.7ZeT;)#0_=SF0\3I=X#1+,TO:0ZXL/HVHHR#Ff\Nb5[@4I:-dU]T#dS
E-&,HRN^fZDAe=61(\F5N-YDO=@0DM-S1)-0^e?)88ZU3A6M\H:AW_76]f=\W49]
.S_T((&8#@J.AY_2K?6[F\TZKR&,RN01MU,&PQ\M(?-+)?5Q1:>FS1B2F82V#JXL
BDOSZBH]<-]T6,A^<-FLdSdcWgB[f<aXIY?2,5P7]IMK#,.__0c#NHeSGKZZ+G[U
f[gYI5Yc0b?L&49Gb0U-68d.V;YIQTZWM??^XaELLSB^E2J0)<:)12Q[BP\^=OED
^H^1OZ>^43eBN(L41L\F]K[O-fRBF<+.fR>9</aQ13Q._^Q/>g0R^7LRJE:L&-(+
MHF7B-WdB_O<S8H>)=\:>.>[+QX-;PSGF.Z/<G:CPMVM8BaL:/V<K/8dc,cU>3aR
>E=3Yf_@[#2@TH?I6Y:RT_RD>X-.5FEM]L-+^ALQUGbGU8,,dB[@4Q2(<L.Y_\@d
3VX#.g+,VeXM(=QGQ0>Y@#VeOg#R7QCBfHZ^FXdWW:6Kd.H0,Ua;7a.P1/dX9//_
LNBa:^D^,G#c[J3XJE3Ae^T:cgPd1VHcSCGK&3g,e>+7^0bH;6:-+Wa3(8Z8<8GP
97[g>6+VT,N0=2>CFK55&->_5ZJa+6EIXRCf_C0\QC[?DY4AKK_AWJ<2X207,1:-
>Hb[>TM)++VQ#;/1e7MPL]5dH)=1U8N+EQ2bC8cND)H6_+&5RUgd&;Qc]P?+_,EA
eT;Q;D1\6/+>WTR?02?4443)@]0[d+McJ659?8J,3DJB>LcdPA-X&TP0ELdab:QI
INV(M5_S-I59D9-JG<W:HS3G)9:eC?gHP3T37>QK]3SEe/16..B0L,T723/96NZD
6(5VSFW9B.-4HODFLO2UW4,5MG?<^<4DN(:(ZeIXeO439LJ.\M,N5N_5P5;E\D:J
cV7;8#^<,5J[TP_OOQG.^B7bP&>BKURc=SS+ME6<()(W&-X?Z8I)Q)S8gSP9M-JZ
KHLLRd^LGWLb6J\)Q0H>]MY9]D<+.Yd1::2YMM11G2LI2KR.L98GZQ;)8WD3I:[,
Ba^SZ[+9Z/^1b&IXJ?G5BaZ\D;4H+8MQaV1XVD3(?YfL.=V032M+B8dUc=>O<+P5
DGWS^.U=aYYVP#6XW;9GU-1:YaKQ6MBRA/8-E+Fc.6=++790LT2HHe.2KMF6H2fU
AbL4S?:2G^?FNXXHeKU5fCS6A\f\59BGIdWP?S[5dEXS;GeKO&&YEe]U=/gSVQL=
]C>>&[(cR[X&XZI2Q=OPK3[1:)d4&F.JG)eLVTG3a)90.F:PW.dYIE(F__7a,]+g
TV)[FJP2D[U\5^(MLHW2,RNRaR6OMUPHc&LO&RTfCZ=S_e05,Eef6,7V3;0_/V=\
(),5QQ<^T]URF7<=+4\N<V;24)Z(Y@_>LDfb2).A.W3ONQ>eeWTACV\A[D#\GJ+8
gCS(6STOXLF,E;GW?Y5PX_+/bT3.?K#:=gb:,,IZ9)QTL]PLZ@ZRFG.YNNZU+a0E
+6=:=@aJF4JfSXOA3&.f,^&d)J2)NId]/RAL>:DR/T@d+F\AI7(^)KPLGf8#eA[Z
#fM[IZ&[Ie:#[M(>QA-Z;1f\c(d>1R@O>AULT0>>aV?/_N9>\_N[&ZXGF9T?UZ@3
3V2I_I5^gc0&b6_&cJ_cN#Tg,MH\<JW#.<gA@cYZ0)f4;eUSLEEJAA&?g,D^&]?O
F.,Q\A[)#]M(R\Yb&B1>GfH2,;8O&7P5Gf4@3=6,^L:23-A2J^+g@>@Gc4ON@M,S
=Be_QHce=/?c71_CEMI6HTB68>G@V=:L72WMH?5/OEe0F45KLTA#(3JEF3&gbR]e
)E#\&?cSKE>Oc]\+]T.A_W,B3I_L,BB=dE[a7+HU9[0GEUH7:Q0FN2=UPY5VR+TD
@BX:T<^A6IOIRLT)U=2Z\M9+/30/46b1Z8\0\P2#,A>(/V>5CVdB+5J7NN)1JAbg
LC<c)PC?ML8]&G-X7O660<@G=TU_M-L?2CA:>ZB:fAJURX+L\S0^E@AO6V?XfGEc
-PT0a&PT8eEM8bK&b63RS]\ZKF6S]cK<Z/g^5?S8bSdg[,@dU6XLK,AN37C4F2)_
1ObD1>ag9J#P-C505:@Z)g)U11;?9SI(L6S6eg#2Z-Ga9:UP.6KV/B#NAB-NbcVS
<>aC(P3ZQPM#^Q\Ga6PVQ?\1HD_AWI/+ACfYO2DM3fZ^SG4(,c<7CXUe1X9dMXM?
<+XJHB7^JQD1=J0Z#1IfST.GbVa#d).a@PG-/+PO)J,b(TF-/dWCF\:Z&5GLW7<E
\>1J16Q(-TU<EP[Z.>f&C@@W=,7UTBB]X>X&AOQ&4CB#cH>1U:QdZ?5=?DS6(PO&
23,RSU2ZW[#:#KUT^N]/J9WQSN@b569.3S[[GR(Q=cd,IF3&?aE#3)DYfe2I5[KG
\?K?ReJUXKKbE0fQ/_?LgZ/3@+#e1M@WQI4IEXD)&JfYI[9Lc.:64E1]d#T2+VLD
@Q(#6OR8LD+PE,1YVWW^]N@+3GRMJ)A;IBK]f1;=@,2E&cY@)5/@QFNP2Z07:9fI
54-U+9PBe^O.eE:<[X4)+X];DPF@De.B1<+_]LAIL3#]/:7M\0OO\1-08@:)XV85
=];F6DNF<Pb5_&.FLGRc=^c?AH[(_;I)2IcJ4@0GVYRXM34=>V[Y&AYB8_?Rd2c3
b;XgWY5\8eQQV7UN5#I&=3G)/UY]?_7._Ee<<;(R@UK/A2J>@:6.IQGO_8TE)#;A
?2HVP4?@a[I<J3gY]O9WKBa2V#(.VC#^<BC@b)Ig)IQg1K.3VE]-gM8Z;65]Gd:K
QICa3-2CTNX+WJ,+BSRU_4](CaE83VHE[MZ#0XO=Y\4<6;UJ\\K[>O3E3TA(=-L+
=D18UNNU^X.MB/1YU\B1B[Pc9C@7dB<BAf:TT215EQ._N57HXAe#6F\DT5J#R?02
_G:eeH7W3WN[=(SI;aF[\;0=P(?-:HL1@HC6a,-\bWQ)X(;IN>:)b\U3]HBXM.,2
ccGPd@,?;\NQV\F/\H)U8IBY\AK)6TeXP=;Y]RCB@(KCU0XUA4cMgP(P:2NXOUc3
O][NPL\Cb)4cZO8(D23C\W+.Xa@C_6JK928S_M(S,71F?AdCd8Tb5#Sb8<>T(KMW
W2[63#Q\Fd2MU0V2X18JMK\?.:V^_BS?C0XI3_,38-6:X:c2W]APUQVDRH2bR3a2
PR7QU<1V7ZJ=MOY91O;3HTF1SX>#^9\;.GI?A3+S#@,-JFUf6V9A:6=dg^_XIE)T
&fa2)db@#RF<ZOIS@aKdfXbSOH66C;[aFJ>dMH-bd[\MZ,I>W911U02GT]-.Qa8>
ec_bQ<a=B4)5A-RNZ<\Y3T/G#[75Ya.4#.GFHP&YA5+4K_Y00XHb>JB[[8ZU;#@>
B0/QdT\JQNDba6Tc&X9=80X7KIYfD91O_[>+G:^B^2TgMZ3;2gM]^[9;0NDWRFZE
(eg7e&F1,I-WNA5P@+O?U<=_;<,&?@E2c?P1,:HQ.\;P&D^g^97SRG0\.\F(H)gX
>+9<8LU\<HB+?_H<f[M6L#A?XIWfLeC-B9]S=\#3GD\D=@)?;(98b5D9=H9=ffgd
HCf1V?0CDC(g-XCOf;L_?J[2:W[6/Q?L\a7/ASQ:9[b#3V8F_3YLE(C;Ia_e9^6Q
<F=S#&=2I@^f#H7aHJU85:O@+FL>QdeWQR/Y8T@@aS3:U[5I2C.IfBca:aPBN:d0
a?P]c6^NX+\<W^H\.H7d9/JB/UFg9b]D.,-YAOKY:Kd_USg(K=(5.699AG&g=+2^
7AJ8U?6@#Q+#4&&/7JEfbHLDB#gJU[JEf;#bR:X<-Pg@7#U75)-@^.Fd7>?:XbO3
&NF7#JQP<ZX3ML.#5G0)dcQ(/<ZJ)_JP):&GC;7HW+&aBD&L-^0Jfa=+_Z0;(;HV
^9HZ]QPDBKdeU+QKf6,=?J<QICDI-c=<I>]C/6d^+XL^-aF#(.K@CcQLK_FZ3&BY
AP&M>#eHY7&1fRLXR#a;IUTC&e;SVFG@a6D:JaU8M1^&551F5\P#;VgU;d.RO_\=
=ID,?SWVdR;@gMB<Kb6(9F]/f9bF\HVCX+,P/^cc9)M-4bK\0G4XcT(/0,4^e+4G
8MdbXQ)46J2=2UF8Q\OSeA?8W?6g)<D)EZSE\ZTg1-\:<f@:J4A5FFK=V@,@13Ud
VK>8DA3^?b1,HX6Y81fKU@3)68;TW>?L-d#>O&b[DeD/?#/;]CQ]A2A^4+Kb)b)^
&HVLc?0aATB[ge.#C)dNF>Df_bP#8-^5dI;;_(d0OCPY#?aRELG1KSaV(:O4=Je)
XEENg?Q=/Q^A14P0@4gLGE,)KdcOg_U6QS5a04=K1PA(MYIHb7JTFe7eCAH_6;D#
e>J<<#(_)?<0TA;@C>)?/2_)?9G[NHSN+Y\;.@@TZ;_8@eU/2gFBJ4;O<c:EN1cA
bgK.54B+/()U;FI;dUJ>G^QK2#VEGF]Jc@]+TZ:>_b_8O)daYFRF1--W+_>_0G#g
)7c:eKZQf7eB+.=<[RgZ)B=K>dc.R?c,NAR5;-MLU2HIMSaRf?GL2^>,c\CGK_:0
AL^GO>8bfG./6EYW2d+U)(2T9eGZJ<5eKcUN\[d&LX#QRV?5BB@?:DY##\JWGMda
8^.bX;:>WN5f;7&;8+8&^:6XQB4UQ]BYQZ0@F]LACXd&L0Y9,8Qde;B1(;#V68SY
7Je_+DO3&/fCaEZ->&D_aOb-QM-B?E([ASS_fWM,7fadM:9ZQCF:L>D644^M/#XG
2_OMKWPYEfNTB306NHcD1bJ\E-cB:-dY;P4E2b:Hg,</K[+EM,NbHCdN\]Q2bK5g
c4;W3Z8OdR-A_Nd)/J1N)U8,QGMXg(MY5BY+LWY,U+dAX5[0OJ;SfbDE^ITURSLJ
.?E4:D&S4b4HG9R#THTR_0WRK+7_291b+=7@bD;\cCE:dfE\P17R]Ge7..0<YI(/
gHW\@IC@:6:5aXMS)8H(-e-bPO8BHAR,ZgVIK@P(04\08.HH,4N-NPEd^;GGVCRS
[BL?@@_J&;Bag;LUf07_CO0W@bLZDLH?OWO,H0T(QaO^(A=I6\H[#6Ng?]Ze=KdP
M,Q>6HA#(e=AT&&9RKIG2Bge3\W#.IFH5e^b[dE?fS,EP14Y]OGdZR1cF1Z55;&^
6-gE&=cdW^6M8S4?fWZd^dV3J&EV437F>E\VCCTA1A((T@/,AA:AGBW70=?XN_^@
RSKM^;0J\L(K@CB>[\1<SW?CAdH6)?@A,7MOJ+/-.,e5M#EI?Jd[^M.>W3(<G()-
@<5N?)Y=4LI?A&bbLTSR4P6FV7dd(7c#?aL2\-M(9F_8DI(P<.&FGS?H^(&3:JTB
3O71,&66X((B+D]S#,C7&Cc\VRWZ8<AR^5^MUFb]Rf7QD@1<LJC0dX5?2??X&P-F
I>&+#QQ)-7.Fd;K.=?<VH8?+BRDE;@VfHHe1N(G/C5?^XUQRBYdK9d8\XDS=->U?
8AeY>X38&_MY_VI_Egd1<[N:E(M56Y/f=f7V:DE<eV-Wc&6.Ge=O=;3b@g,K_IU6
@>]7P0YYaXL@UO5VD[2COH2fWJ@39+J<8&ONIMga0AA;2YVAR<3EI0FLN1#S^HJV
W+D=d?8H.(ddHQBR?-N^&@/@_MYS7FfVUM4#=3gU)Z3\gFCOPWH.b?Ve@.?DJ5X2
7;E.J4TUX^?]0eD1BT/f(AEQ=TXa9b02g,.]_7K79EW5Sa(_0[T02I_XCeLC)0G<
+<?2YW+P1^&].JO1gg?1-1\eHLeAJ#=WN;gR9J_=a;\MOC<5Kg(:^aGab@I1K9]N
QMg-@D28GO#O]/7O>G46>AK1c,J7VdcWa-+^.>/c\:YF?X<I(0JK&D#V4\RD[B?D
L9=4D#c@7->;ZMCVX/PVcANW-A-B?fF-d8^27b9B;^Rc,e>Tfa@8Q<E39\c(aU]I
7&3.#105U:.4Wc4I_MGg(;239I7,Z.2DOfRWQ?L15B>aGF8NDDG368]af.5?\2]6
CD44Z-c/NYJ8CdaP3J7WM<S<4e7@-a4U@7DAfdTR4@56_(@<Y;RDM22T[e)-N,]8
b2&^I<<&RMH\8?<:V-VEXW67\2<b:TE#>S+I<4e4\65ILMOS14^:HAf[KF8<fg70
YU_CLG]\+-3,gF)?.])_]SW2SVO<F:@0f8037;8@178YGDQ9g:GXPO[0XDI[OMM>
CW>ASgRA>KU9H9@IAdNPdCM.3eT])R&GJ2F4Kf9dB(.Fa8SIT1fcI@-TRQLbb@fd
Oaf;_;G]_WAH[X,2LJ4[H)1DMd9E6HAgf-5/HM#IeEKBRcJU5TX][0eF-:^/TCg+
^13^RE1M=:J-.)e2fW0)7adT([II?F_fDHFL\F_ELF6;\EDFGNK\3f=,Q#(G5Qbc
?R)CBWd-##7;5I[;4FA4:@GJ8O/\4@&Q+<XN]2^CH\>)RBZ8DM-N1IPCdJ.8P9TQ
B4a\#F0aB#CDX;>f>WeB2VA+Xa0X((M1Z>aN2FL5,cJd^CF^NbDLDd2DGAYQc.;@
2:SL22FG8bJM<2GR[Z96KD[<_,LWE(JGC6d8TWC06,F4@QUOV2e)5&7G]BVHd&X6
U(^_L#];ac^dI]:0d/#b;XEO13L8E7&N0>D1-bN7J1aFX+\U=X^J_HM.?2P^-8g6
)F;aYR@4+)&<?\g?F^]M5P]3gPU,+Y29I-XCV#D-&WVQSV:;/0PR84;LL4J:7(9+
A6P12/3f_G(R0@dg&F6)L4D#b4(e.a4=ZI(E?e\MGS6ZPL>+VB2A?2;?&CJb6JZB
A,PcOPTDJ9YVJ5V2>8,_(V1bB2B<G//W2@=/^dF[]IS(E\TC2.,UP@dICNa(_B/D
3=6)(:DGPB#+I^)F8U1375Ud^KHDgdc2S]TXC]#DZ]EcD7aU/dcYRHO7F-Q@Ta.R
2-2EUc7>d\Eb.3N,bWeaWWT0?_Y48[BVUU7KA&/.@EageEL@HS(]ZGbdM-GK5PGU
C,8&Af)\&eUSA>=HDZ=e62_dE#fQF6U^FI0.;[fc:QU[]\CL@>^A37&>b[&AM5<R
X>YK)=@5:F10f,NX]egYH^I,R-T>^.1RSIT\P-bEGP9M^U)O:MM4(R50OX?[JZLL
g?=E)N3?EQfQe#S70B\>EbE;#XOYMK+L3\^P,PQf4(g=T<;gQ5B/KW>-E\S9Q?SC
+<B;8AFX)V4U8]LGH2Z0/IJ0M<.M.=XG@51Mc2G#[MWgV,LT;UV1?\[6SLe6W-bM
]I&5ff/;-@Bb+9C\M<?AV\?(6.C7Z2R?KVb]BCL7W&N#MY)9VZ6B0gOTR]NBVNe0
43LB;6+b@9U;/S\M4]<I+d>@,7V]XKE:5JC#e7PK6M^25WXg8<;EFgXP@ELG[Zd4
cG@W(6(Q_Q6;D^IAgA^#gHERE&\YCPBM1b,\NU1#:GE,RX8bRF(71SMfVWGO_>+,
e_<RQC4Z]:P(BX9=Rd7D8X@d&.SN1b:Xb6>FQ&.eK)0F/?K7CM_-SR_:Kce2_7f2
JF49^\W/WaRB1WfBP9=6_9+&3=.O-N&c0\XUUMCW8AM>[RcGNfZ&bRZf]NMXJF>S
Z63_d>33Z=Bb&feP:.+^T^+S3VKcc4;da0ePH8OMaM2.Lb8X3#/AbZA)KR2-b5^G
.-HA9LZM9fJ],ed<e8)e8Zf-82,>0,F^gR&X?..BJIg1M8]eb][FQ/E@WF]XY(KF
2b]R,S\JY>QWDF^=CeD/^47[;]0<@DS5;OZa(&680HEZE0C+J:I5c7A]U>GM+X=D
NYG\[-DVOP:XeJC5UIDWc,V#).=#S;8^O.YE8V0<&;D\0VP6=4V>#(YUFCT;PULC
D:LMYd-=RT2<<R:c9Fd05ggZ8M(Y^f.Ig7XeD-@(0CNTdB^7(5;84SNb\Ca_+bQ0
(>e-,C<&94;]]D[<(M#\eg;]JI#&J5[KF#H;]/M7,O7b_FM;Eb,A56A:0PAN2AUe
bX4FCHY6f4LGbVAMCCE,-RJK]?BQC+CZK.XS2)]+Ze-ES\IKgO87Bb><A-H7gYab
:9\X.F]A/3=Z]2J-8(f2O3^[@cE_9;?O@N2OeF.@SYY6G^XK62/VdQBZ&5_AMGFK
#fE?DE2_8LO6EZR/S.WGDfIK8Bg_a/c_XM=#V=]0(0;-#N_C3,1:+R4Rc&f)^C@X
G@\7cg.K?fJ06[EV3^FR8dJS<8J(ZPbP+E8QX;L(XY?2F(+&M)?XVfc#b1/ZCUF:
?XQH31A+TYR578PTJb)&ZSS>HCW7-GOZRg+a1S+LWO291YC3Jb9S>(4TRR&<dN_=
@:5Ma3[dZ+>(#4XV>JJ2e&3f^MS/_,6LG[,D,BJb4I;O5QQVHOUK3(\\E)P&)GFb
MM5DN@#VeB6@QA8V<GM(7f##<6K05bB>9QCHbQZ<fJdgA?=0;,RD]a^FdG/@7FI[
aeaODD6O07#;<57<FF&a#0^:1>(9)C>845H@XL=MfZB(.M&d=7Z.+GOE^/U-1g#D
]=U5NJcP-a/RAe.#KAC[]JcI-#7PGNbS)Kg^a9D_4(b_PW6eCU-,P,Zg5>\e2_>R
f&6)Sg83-;IQ08Z1Dc2SZaL6c6/87/8;F\>VW:3/72Pb3O?XI\>bQ;OJ#cbR0fZA
AB._P2GWWZA8G/\;A[?H5YIGb#6)1^=QG.<c>F6E,/]LJC)cGLcV+c[[Sa5Ga,](
BW&Y^AY3XK9d@\cOP)@L,?UU\\d?;UJb2)#38;e:ABJ7G?Y(;&[NIZd;JeWde=PX
I9HR.)e-NZdKUR&BX8gD=NC?P4RI#1PWA9>O;0B95YgJ2bXf-OJBJIAGE)_R1a2:
d2+CE=G3VXH:_2gF9=(O\649^=7YfK=5LAH3eQ4DWC9=YgD2=^UdC6S-S1f6)NAg
@@>4^ZI?]WDE\#./UI>;=C6<ge.bgG?M->3ET,:+5a6g8Uc(\gYEeYJQd^Pg;H(N
ad=@<]V/8289@<]#9RfID6AN)VH#&;f7X[/B7]aW^Vg&K&CQKV:Q?F\F[G\)RHR=
+0]Pa.c<faOK9V#1]MDP3U#?91b[7-8YZB@W]]+9X,XT1BKI?MN2YX0QVT^Ac7\Q
\E92TZZR/bPO74<@\3<EY,bYf^@H;;/6DYI<TH:9R(RY;&FDP-+4T[FS,8bLO_]C
ZQNQ[Dg@g\(E&GP>V=4e,<2BT\Z_ZTeTB=7EgIX^Z6f8V?-La1(P<ZJ>4IX#WCAH
97J.]IC(P3EN[DfSY3LG[5cf8aVfHf^_KMHFPe48Y;A91fX7<(B1&&e,3#@0M0,c
FCV4[.N1c3Y?Ge=C38#GD]157FXM>JQ;8f>#c)[/UWJf?]7\.+JbdO?UMRW8#,-2
DLSBE<0Ga#YD^J1FYRZ557,O:W))8NAU>&FQ_c0\G9H:O:A+AAD^Of,L[5gPO+_R
7c;U>3?+CH<W&H,K.5Y0CN5UY>VeA.2Y;O+<2MN2aBHFNZ4P4V&5+bDFe?+#INMS
8+A\G)GYJVJAQEWV7E.OD))\PV/2C&1RBU#9(H-d(<TcO0VFN<.(E#^M.SS8(<7L
[Ua-WE9&NWg2N0ZIDI]2IS_LO5^OA-J3<e6Hd7V]UZPWd=:WSE4P;>-/D7(TJ1#9
,QE(>]UN/=,>S\Fc(>-.)0J8HERPEW=DX(27Y\L1CR9+/B:\ZAc7TXFPf<\)TA[/
G3S#faJ;RFWY_9Z_/Q37?<MH@d</DA^(4GG>X5+dUV[/d=QD4SYfO2S;CQQ:L.Ga
#Y\L3aIA1.gTKZ7:1_M.aZ/BTI5U9P@92.>gVcIg._FJ@beVBg1cJS#[\?)BR_;Q
>+gFE9J.9@;#912^LeH40A)JY[=d.9+)8UgbBPg)U6BX^-cL4:[geMBO3.UZ/A>\
0/?BR;&5B79E=<SgW+cc)J.259^,9fd>8]\<E#BR#5Yc2Y4gR^O\WSE/]::B.RQY
0;?+05b1+SS/-=JFc?0,_1)3aOW.&?W=R0[0g.9WZE,[3T&?BObNWfK_2Y.e2#9@
S0O8U@Q6e9FXZ>=MgS[dY[M]T/&:<0A>#2)VV\fB:1MU+Vd]V>QC<@XEMWL]2bH4
WOb(cZ429.+_^3H=C&]c=@R3^YHa;35@Hf\KgfVL1[#@38W_E^9gTGc5#I:&7S+9
J54:V)>QL9(HJ:R1Y8LA8bJ.10,@7X/fde/[b>74A,.1Fa#c\T06Qb6E.Z7:V<M@
QO#(caEfGIcT=Z[#N[><_0fecS4&?@Ubc?SW@eSFL[#>;>8G#-#1]0QN2N)gbG0<
ERM6cR-UcBWL@6Y1-/?Sf&C6c9_YM@=+K7.[+c:YT\Y#73eS4c=;><3\B\74R))G
9aC,XA9E7-gRd6Q_Md_eOGZWE19B(T(X-JEcH+]Q+,<;4DRB&#KVE5[5IJXa6C=/
>4J#c(2?Kg8^BNCT7a&IBUHUK89]3FV@28W7=NU(5B4UN,b,3JK,HB=YeX:YLR3N
-c:L6405VgYQ87#@#9#L1_MQWVR.8FX_?Z+_d0-319cYR1Wa)5VQ1)PC6MK4-7WQ
J.=gg+ZQ#K(6[G8XQGD(AM;b4>-+X-#TG_G[:C1HcS;AT00&M^9=T]Q0\U+_#-5D
31V9RE0IQWZ>JJ]L,U+]B]Q/.&b3Z,<-5CVF0O8OVdaRQ+5Hd[HEJGJ,B_Ze)_aJ
Q,=cALT@NPN:Q2W#DeU@6Kcdd-T=bQ?+JDf650(UNO=-N6W>N5E;^.59+HfP(>=K
&PL^gT>-SdMYQC8F7^OAH=D\:\.&O@D^HIGd2/cgP?g=IEg)M9I\2L/DO)CG=7;2
,[Sc=4dHE]G3V?>dI8fgR2ST?;U:J[[LL2(aA;,C[b&/:.aDC#2)fc?2BZKHN27-
3g\1gM#R2D)e^<HW)d4LLZGR#P]V9dO;a_#TJ<a&W.Ac#Z.#EBN?>8?CV6+@fgH(
8+>DWSe[S-O#8KYNGY]R)#?P)89YPf/1YDc=#/;+9LUL01\(-^b-MN7T+A&1O>Lg
]_\PcFY^U8A=<gBXFZcEX&XP17BA9/8\8O1-BOc3HL92DWd9C[ZU]V\IFGBB1WP3
a+K02.D6I_])Y_[++IY;GgBA)S9+HT\FT#A)6.ZK8H<A_+0c#^f)069AMO#?8#)>
:VA)V6fAaWbg4(7893X0WJ0FB0&,KXPU;bKc^YAV>W@d)80FLQb+;QJf2.f7e4#I
Z(><V5V9]6>4a5DZV7NVMLA3MZ=28@:(5HB+?B[^(VC+g41X+L[DX.J-SLMXE_44
C<XNg^6+e0?M_U>d41C?98PW6SZ4Z,cHV<)]CX.Me1e>LfSZdQ#^=H5Ad&_E[KU\
IT4dJIU[294KX@39&KX1INZP?b-eVb8OT0OIW;+aRZbgW),0I_V9)\;;NWAE2S>c
U6;eLN9JP7YAHWS#\G(Lb93.?Ag6?EO4KRB1[c0]GN@Fe&Xe1U4RBZBd[[_&e^\@
P@#HeQa>E[<?(4aS4cFW.^UL:W3c@aVD#,:L]M6_cD:#(V59O]8N,J(@LG/E7c/:
.G\bc=d/_b_DLUPgT^U+db82b.2^46Kg.b:4#O4aRN]XHbG8HU=_44F8(AZ[1db=
Ld)KJ=LAMSFLF^6D<_L5/?WHK?1G?5dL=:+gK=[5?9c#PA;T(F5(AS0BY8FB9Y/1
33Y1]U(e-WQ;CSJ(bYJeUda((4e4cZ.;,=KBK.3&,dG1B4/K=gJU/gDAO5;B)JL?
)g+(b=-[DK3Og81G.[=_;G08XBMgG;Waf)7Z\OaEW_#C5^cd=>4/<__A.9<OBE6Z
WG\^U+cE)H&P4@:MY12bc2QOZ#NO:]P.J<5cN9G8U/g&efB10(I_[18)<+(<0,<Q
7EOSA^e;)0P1+2SD,7MR=4=KLe-TCD-D154PD3/_c0-566^?DW7<G.?VP7;OK)^c
8UD-Y]QJC1W#cNX5Rg[\g(:Be@;4G5,U?0[E])_Le8M3Ve0D_L[,F-P3-BE;ELQf
GI^5UP3MA1HQ)2>5Q4T)1+;aDT,([VFK+9=-2@M<21@9XTd)-WDAJK^9VBOP2;HG
^>&;e()<3]?^<^3-\>K\1...@P1OSgRZR)VB#fc:4QcU\C-7SRdcYc4]Ne]fTT^a
S^Q;\2aF.0])M1]<HN9=Vced&YIB+-L>/C2BQ43VTJ@)8)>(XMfS@SdUP)Ue&eCG
CI,GQQ>9)KN@6N8XbXB-=>]fGaUW]T/g3UI)&I=-_3DR0F=\I8UYBeLG@I+2WJ,6
WGIDWK9.(_Dc)JVBea=.3c,WBH@E\[N:202MONLgN=.P\],1\7;1/Ng&0L5,NJI(
8\K3)X0B<)bdSSPZ>20?H6-1Jcc;--=g,+#TZJMLX+f>Wg;XBaJ-K0bg/)/=#4V7
Mf^/X:MUJFc,@C)c1C14,PW2LQ18CO><-_Ba\[g_TC[6d1]<XZ5<SL_S-=+]G>EB
J-F[M#2<6b3^4ZBRBe7+-,W9dO(D@59LKfB2,VQ\IEELD_Z-TZ8:;EFRL3^V_baM
;CJG+B]a>^-[]MJV&[ac6Q#4C^QTaN@1XJJMa,^[_Q9_^HC@>bHYB(PHJ8A\8\Ba
LQBLZE)c.-XedL;@ZG2M3;;M+B/L^ce4<WLfeP]&#S/@N9HgE0]E5/aa;@PeAXU,
Ic7UNN\g]9gEf#/WUPRYN1A4,4#a^,GK@7B2U?@X_&W@gH1O&7^28D@A+W2FJBc-
S>1d3O(7GOQKN>IYcPO8.Q0ZVOV?a80.K2-6((&(AT^W>O-28O92TFJ]A=PcFVWV
Q)2.9bN[+<>^F?NL^N&HTD^K/&#f^E9M+\[ccYd)N;7)2W\7f<9Z;)/KV]Y1V.5P
IXL^W-W10f[JW>d]SBR[U5C,BR1fIWCE5<d3d8e_V&B@K40(BgUaF4I,I92^]54d
0KF]f][2F6\3D-5F;/),bUV#c_5bO(0<NTcERB\#@)BS+^PFad(9GU#Z)9WbdPC5
G5HRX=?:)LDbf1@2I[/+-VZ#T4[2\3?(2\Ia??R#&DMNN(cLO^>=Pf5g<RN.gNBb
VHS\T>_K^@AgLgaf8E]M7,)f<3MecB.3]W4PRPKGCE81a3-)RgXb:03-\:-O^)+/
_VT/K-]2DBQ3#8,&JLA3<B-4Q[I/#K1]9RTX72MS_H;;61G..JCX\5=C.aM2@XKN
KX8#IZ,aJ=/O\8OaM:(/V39]c6NAb5HF\1:Gb@dWb64L)W=Z:IeKCVce8PbDPEK6
e<2a@8(R/RagK]0BQ[dJFf\Z<0ASH=+WXQ-WT4dQ-7OMO<ML:@]g#6Ac&]BM/Q7#
AcLf^JV7D\\FB.>RM\Jb3FH_K#;,S5BN+bB)-OG,NZZb>^0^F_--WcWA153a:74F
HFUUaAeWX.f>TMgSe[e8A9I[1&eJ#?_4)88K6&L5-#b#[YR<OJ26SCR=ONT5(LAL
e+O#<@-.PE\-W2[UY1AN<g<XPdRC-ASQLRBT6&T4=/V;\/^LW@cHO&XOED[4>:M>
8JNF/;,XTf)E2E.->-)4A_5V98&XRe3Za+_bb_Ze./;E7F,I@AS1X#g7H7RY?-?/
eY\Nb6@=QK&I-N2NXET8B)@11Sf5Id_8>K(C8\5GGLR\T5N:c^gNLNHdYJ:@4bW0
C38c/IbU/2aY3PG.YB\4:MI),?Q+JAZNYA_Q3S\02#(WcJR5XMb2-ZEA-YREU9-1
ae7@UOL/<VC=-FX#DH1G8CN&?SU0M()LfCSadU1;&9=H1.MNc6DP#3^[6TaOR0fc
4<:3CO-5J96R9:_A0\.3QDFLUXGS08ST>[HdB(->VS,Y?bPGU.HNLF]+9.:_&X0P
CM.6a:&_OaSE:1[cOcGc56M.H5R?MR(+S(+QFK;@3De^B9gCe0/LEF/U\-B/[cGc
TF7HdV+Q[ZI.(dVMeS6UR7f0d:3S<J2S;6a&9WP8E&RZI-/0<@NPA:=:K5dTWOST
D7Q3&_6HbXW/L/#[@T^Pb4c,MP:N,)]?#]#@T/3<?+=E<F4W;R.Z@_;g=]#&.7-1
[>Y:)aeTAG.fHPJ^:HPaS8^TMOGD_cWPY<DQM3-0^O@P>E5GR&PAaI6;5Qf[B)5[
#9?f<=e+fZ;YI\dB<b(4J7G=.:E/][EHBWQ#&G@A.:D=BF^_8YY9J(_66_c+>gX=
[U<(^HQ[2YGDa@]3_3WXe@2eZ2,K,G3:#>Qa8Q.cFW66P/9AIX1#7ISX5GN</K65
N359+B_90Te58#WA)\BEA]ROW0V:@1e[IJR&+U\E[M2a(<)7(XI0<9cS7?\1^=JM
^\.G3/?_=d;PfPc,EZ;(I6=BfAX(^U+M_1IU3<=O\(ALQ7Y(^Q)3-J-eAUHDaOB2
K^0YWA;Q21LW9>d\0P;CZgTFOb3D(OA,@A99-P\f>)-X.7,E)?,-1RfV>RYR0e]T
UT=8Aa^@6,)2Y@MKS\caEEBW9O<E;APY.4[gaHQdGH//aUG/L&MM5IZLQQgR5XVT
&:M-+0RV^ZI@fJ.DULM?_:X6I\bK6+4,H;[d.Ugb<^GP5dUeJ.KP@GCG]0QJ9a:P
47]4ee+BGIQ<-6\]7M->?KVB-1YB\PQ@]Z:O5W@NF:afP+Ifc>KUOFV__R1^#^c1
-K1@,QB^(2Vc2g8RG.(CN2G:2J6G>\\F+-4E^-+)2D[,,N,GUP26D&<]eY?N_AT(
(Vg3d#3JbMAQ/3QAKP<(V:4^EB?YI[@GP:0ZWZ/c^&bY[9f.6Ac[=bDdY@+\6MC)
@(>5^^IW\#BBVgD<1A[8\W18\=g\_N4<:DYd]&S2;>7_LJ:&;N9RAH<]]33ZQ-@R
8(]9BHECL;H]_6[0QeU.fLZ,ZW3KH><QeOPf8^e,DdM5#P;O(8:bG+/\E#9W?&aY
=G>eRa-GDe<&_3UE@-([&dP#/Y?Q9U374FT=c)E97LfU5_1RC?I43HL8K+aS:=D1
JFW7KJY3g77C3>RYGA)UVIc6B-AYJZ&^VITfBdQHg2V+;2Vc(]2T45bR>+6AQ?-#
Q\-QEW=]NV:-SNTL51#_dHESdRLTAFc[=5<F5BJ)P@D?5]6@GR[N6FAcB6@:^V5?
756?e+O-2c)e?T,)gfIRU@G,D7NWZ1^AAf@S^PO:NDG&_G8GWR5-^=YANGd[N(7\
3gU6TLS.:]72)<_DYNSB6O):?A4JKGfT9^>Y^U@(:VI65NgZU]0<PR_H>Z:U;_<7
XXCf.aU0B>+/RG:\OJa3HY&3g>dCVa=#=g4)9(^<&:?JFOC0@M=UE3T4T7E\UIc+
A_d96R6PbG;Pf;e3?@c;B2Ia9bC.I>-@J45Ng/e]d&@#bdg6.MN/12#eG<Q<b(;7
^[.YMUO-&b8:2VSJ;gQH7fHDZe30[=(Y_8N::\_daeX58D#X;NeB.FB&P&_Q#-cb
-4CB8f,6)AY]2I;=AD2dBA&M[_=a5&\#7UF3_b&D0?>TA\:ZIZMa#_1VQU5c&2c<
ANQ27A]_/a7T@4B&W04gg#/X5GN74SS0W^d3[HCI>2:IQHBI99/>#1:;1<R1P=AJ
9@Rd.RcUc\;<4b?LX@O:1V)^6CD\1B[GeCa=\N?(VE)G-=>-<2&[>c?FcTg(&Va:
W:B\R#ZcR>?XTO;gK/CgROLd=EUHC/aYBR=O-V=9AOKaTg,BQg=2ba-Z7f/Y0KEa
ZSZH/1>5fd.?cTFM>gS?92+7&Y#)>AeeQcHF0X(,=WGQ(61:49-=gGX,aKSO^J+C
d<LBY^(PCCGLOYZ-DQEd#N(T?H=05QQ<W,&]c?X_=Y7N,MOG4-BfF,UaSJOS5)D>
:79D173OSf=IdKXRYAeFS56)5Y;d1H?Y^F.JS>]KGQZZ&R4J&2,2Gd8ZMZDT2F;1
JD2&4.Id\/@0@V0?9/Q[B-1R^[JBDETJ[RGO#CN_CU)(IQdH/7d84JXA]Xf1EXYV
/Wd^<6V)ST2cP<H6A9C]HMXQUJ0X]-Ee>@_J3^_;(IW]6N(^)Ydb[EU3&-<]<G6]
9U]gI_>Cdf)YTKXH,c?7,bB&[A#VCA6RB2DH3VG=a_3PTE6DEVETdR8NSf&f4]g9
D=Ta56HQd7=c->N_:^3.F#f/-b1JAWZA8?6W\8SJ?Q\\R=@F]WS[]c=K\H2R,>5F
RaI)JKMLVF;&^6EYeB#cNQ4W:.0DK=6L>4dU5V6::ZA03ZL\U-IVB-)HNfgEKe+S
b(K)7)Z&D#BUHPf((6gBWWV0C]LE;IBC\,^Ta)9Jb/^17&0CVZ-d?O.K1b8Ob^GC
AI4&K?SJIgb96)6#A<T5C[J,NR,664HG/Q30]aRDV_(FH?+bca>/\C;fP(C1<0dU
eVQ0I<T->@&9SDgVA+5OeSZG=.)(7H^BW6TIWDM1HdgVZU&849dC]=QgFggQCVSH
T(KVgTT.;((HM>ZBC]#DLV0XLWLB^T4gP[EM37E?LA?)MWaETSV1KTa#FKB?H)=I
;LRS>Q:(P@#cF^gC59/5\dY:.Jf4AO=.Pc>OS6=S_e5-7_QbRc<UQ&E5^8Z>ZPWF
?X?4<.<TJb,Ta62P^JC9/2;N>00D)RI;,8^a):,\GTOc/:g3WL1dd=GO1-N70&)J
5AA[SK<<(J_Pc&cPadVL>T0XFQUaX.>QCVXF(Y5;ZJQXHT?+ZD0S8=7;)a(c_Ya2
TIM4Rfa_I>J+9&B3QY\aN1)fANG:L#afRb3gD,)+GFIEVG@T;G4X6RKOD,b_MdI2
fYg;EEaR2YS06-^dT=]c\VA1CdE((@J88?WF-Z>LU(fO#21JYWH\?4bW61WH-YH4
U/]U[8[(1If#d-BP0;G],<bd9U-S\aK:S3V-F=<MLeT2>d&^2V+\T7,54aNSQ#)S
0Mf?K;fGA)=^d#=Ib;<N6Z<O.JPf(YcZLBP4-ZRDc:g(G.F]Se(K[:&0\g5#[N,G
VB1FE?-92fR3@T0H]dJK9(K<_^-U66HVG&Vf+:(8R)BZ4_\4FWS-=R^JUA8]f;^[
g:F9-J;_dXDZ?9FgS@MUa<R6ET9U>?4W@\:_@IUQT<+EI[]4bS22=W[[eG->?#6-
-\a2c-4>/0/MQ(^C8LKaE?>#]-:94c=D5RZR9SbRY<K9JWbg849-D10ad4bN)=9(
1+A.:.03fK9c>FK>F1A.+LN<>5_XE>f:(UZ>7(_NOJaBFegT4T]S;b:6AYXLJVQc
<W\KRLHO#?gYbEJARK411[d\50_@A],0O]Cb=5]@:PJ)c_EKb[6TJ>IX8g6a\]9b
X@4)OTLaZg]NS,>5UE^+A&&_.+H,6/#WYK&_-^MAMKJ??<A_)R;VFJTE)7/V71L3
FdQEJZ5[g7cB/8(fUd5g9G261:X1PIB@F1eZQeTVSDX&SRW>1UXUbf,[++MT=3J\
7T<W2KH(_fM);gSR5&=+R@EYdg#/T]+#&M.]G<I)&\QV&I/49^\]BE1GXA()bA9M
e15-\5TXWO_(dIEL\HI=R4?5\1Id>cYUQ0#665)c7eD]6A3B>Q>O5QSE_T^]FSPX
Je=KfINZ&^=Ece>&UG+-G^a@:c(Ug//@8,6b19S.75\F,,\F_/eVLeI6P/5JGY.(
Z1,7K[LF.ccXfa_^eQ7AW=BcCY/:_P84=/G.][;7VCII/?&P>.GcURaRD6E?J07\
<^6B]B2K_>H,V8P-L[bLVa&^-<Ncf)_8f^R=6bVDab/JG34,51;?RaTYY99D\ENM
[dG2A<GV\&<:NS]?EO>@9:VfPPOO=2Pec@Z5/\##?U@8IME2[[3]<0D>3I[=G@\M
XJ+>TO;b]A1Ug&T@WRL-1a;R#IT7RV(M48XHf;Kd8)2+4dRF:/gJ3aXB^a.\(1E&
Z),dE&.B\Z-C;WQeb^VQM#g(Ag&NY>D?D=:fAUE:a>fP[H^E+cPg_KMC_@05/d4^
g6L@H4KYf)F:68/O9(Af0O#ML_2^cceN9XFEYS<O]FX>7abL.1]5\YPN&bf_fOL9
VIgLa_)c:G(00Q:C0aE@^X7#+:GOHK=,SLV-GdJe>Ed@5[W;1=9FIQ4F0:H7PTdZ
?D\d,_.E^&K.fYHR:I-Sc;K;06D5&(I&dI_7[BbM=cf:?43Y+TL5@gYL382--f6Q
6R1R8=QA/B^DG3)ZB2DUgfTSZ)NVWF:L[F>aBIBLa-+20-X\?8\W&G?/dH9b7T6E
gI?3O;d^V]WIQPZFQH&GVYKJBE?2#BBY,d#KX\a@MKMf1/Q=Td?_T4^<QY\+K[=(
&0=6&?+QbUJNY8>Q>+M3MD+A)XNES[)RW<WYM/5X-I93a,M)C32<1;>ALC;<_OR+
A]Q;c57RXcAQ&TMBDYX\N4_YR;7dc-LGZX2Ff0g&+2^fU6]RR#K2KF@K;;02Y0L2
[R>Z]NUKd_<4Q0-bGE5(7a<N9/U:)D66?.>G;6]U1ILF&LCXWAKRCc1@NcC7fdHF
1IU+f/-GU,Z]+3X)P3VDJR;1]g0L=VdK=ADIRC]>:KNK8N&0LIGcA+b/6_7YIZA]
DF?/g/G,H\^]fRfHT09[-e;Zd,A79D@+;,VFCCXFK#751M(MPZ^T=W05AEQ3_1\b
NB2c/E1I[^CMb./O,J[7]V[2^]QO4&De<ME,#\S[<B,b[?&YKeHcE10dC/189):Z
58+Ca_]@[0X,U?eaROLW\D9R7TGIS)-egbHO;5&^X#7I^bf4ZGWQFeC_cFL6E-[K
9Wb-c]BXRbP@I\<.VeBN_:=1,Q(E=e<HT.gf+_WT_E6)A50c3W4c^AIcDV@1OY<b
I8g_(\cKQcFF6=E.)Lb]bcJ2,&4M/=Cg]#2GUC(BANQQ08AEMe)Se;0D_3cG7#GE
C&bg>&dZWGg>dZ>E#]H<2QY)[BKN#7;Qb)EfF;454cDZeH5Fdc/F2O.bTF.:/R9Z
L4VU<UD<[NMRU8O9]2Fecf(M6TL(dAf7X:(KL,]GbG)J88-5W0M^?BR&1OeJg1V:
f-/@UBc8f(L=-c==^4MT72\K+36EP06d\23_JUbD_9KI7HPA_&EKQ<HF6ED79@#)
ec(N?KT2;QH62L1.OIU=]RCYa/f\eLTM)/-6<&-:F1fB;,AC-9^O)cE.OWD#Mf-f
Ad_E-,R8ZEZ@TgLGf:57]Pb)4?G+W@a/1K(.D>T7E<>&^US,(P3NFd\0VA?9gB6[
aPWZFR=P4MESH&/9EE;)IPg9L041#01GV(@,e4c>/9VRZFfR].NeT]E?-LI(C(BJ
f@S,?CCH8+@XCe7B7-DCPV\W0WaH94g0QVH)MAUFC3d/E=)MZV,#M)gWHa&2=.<(
,;e,RJ/.U;F;_c)P^[8,;g5De1PFe5Nd+YJe\CJZG7S\>YD38ge;[=U9+M0@fJ8,
W(d,QGC^)=]BW<IK?Ae/Gg=?4fO3+4c?1=33C4-S<W]#>2FJ&eX;8XY_>bQB5de>
YS[X1;_\@:QC2bAW8Y)CKLB5E;;:)?K,7E>K)[5,<cKJD?2FSDETZ?TJ:2?CZ\00
1g6-VCBdd8P0&OUK<FY5b_T_>#e9KWQ9F1XVY8XfZTDZYbgOXV(0<cK(@=T,@XT8
CSO4Qc1;eD_<fYHDB8#\#@,dX9:?ZLE8W\HD0JNSIH((4LEXG;^.HAS(KR&V60DW
Y(87KEM>c5R?d\f,L7EYS+ZU&8I9TdEN2ZX?&>[\B;I[^[&N5__VO1M=d4#+g5[=
T=3X?^?0=HTgdCC1U&PKZF<\RTc/,S(TeE<[=e.2XOC3=QA0,<I&MLJUc53-H.5[
RHLg;XD8]2_)D7&(U>7O<CS@]SS;Q^/BE?#UaIZ8G=XZK-D<[fDRLV#>\fKF+:/;
F57K\D)9#ARGPUJH3Z?0AHe4JUgd_DI:+>RDZd,?J?HJO/._c;XSPAN]-ReM6:>e
XF?df3[C#W^feS-&2=eIZU/^4V.UIA^9_>ZQQ>917U+/cE.(d]D6+Kd;Hf-I(],D
aV7[03Pb]d^U44dS.1#:dWMKXaL.0]LP&<+_8V,8e<M[=J.@>]+3cQ+>#J-5UUe#
eP^QVZg?SgXOK?.VI=W=8HU70@F38gO73FN=(AI(A\\>(FE2HbdHK34J-[0[TUXI
6&IH(R990G>^1I#_H>L8PBa+G]3:Oa0-E.e\W&U]5@VRa&N<GJQV+_=N+RW6FA.,
Z>SVR^/(FD[OXO/(5MF3H(DB52N,BU9B1:395NAD4#B1-Y&U589VUTJD]2IC+c9N
1JeMe_X+OU6faT+N=)N71:V\cR-X20XT_a8]\\eM?.(H[YROK5VI@RbRB[Ne7G?[
JI@KSgL>G7KEC:5bO>XZQ),gG:Bf?G.PFI.D-NO&@-f<[cH8>M#WR2N1)QP&A=+L
I_]I00.KBXKO-2=>^#&Q0cN/[W5R6)9=Z&W&_6/4A_94JQ-8cF_Z:#\H)\ZGD7]S
#Z?1:fe\.V/=7/E+-(\&#9+<:S[A:)d6TR^?R,QXI/N_a46^Qb?G2f,W<7N.NX(Y
-49/>Q?d&.J&9@GS._T/c?>MFA=9gBQeGeUW#,Ae3H8LDDK50(=@E[=e>6B+^Vf_
f./^T5Q30W<#IMcHeM4Yb7R@bgbLGB4(B2[<)-@)9@IO_c=WU[857CS<XWIcY+De
@R?)f@Gd+1cG<&^cWZ#)\]GF3BZ_(:I4VF&A3UZ(THI]-5,cC(AJaZ=;Z=GVU-6Y
V04HOZe4ABH4:^QMB#f19RLV]_?RKFN(4ZUa4,]f4\46R\>e^BP(K6684CQ8XfR7
<,@:282979<Kc3B8AM,;#TD<US8<9P1),b<fHRddY15K.cAg6>5UO&+)VI\fVBNS
Y(N&#/MP8cD)EK[:<2Z_:2B#8:B/48de9_UD<UA[/=;aP?F>N)MLO/_6\Yf\;=:J
JFU50_;^02^=UNgb0:3A;KKfc8\#XZAJb)Icf?L0\]b19F9HYg3#W@SH@Z;F]H&?
)5g)WJ0=a7e0gGS0gYB_L(-=A25X5R<IEdNIg=VB#KGfJG;F@^CJ=X,77]TcLdNN
8\<+>=&g@ES>_G@C-<AV]-?J22<(:=eMIN)B2\5Q<5&5^\APC32eI>_aMg>^#=bA
S94/A&I5[KBODG54D-)0_<S8Wb&HB689^g26=LAc@^\_HfdGMF_DLS&@+[EM9bU]
g4K8W5,ZbH.73--5B@c>)g=<eg?]XN2FCPUA,c(LA_e+Y/+;(bF-,YL;GOPRWcXM
I]K9,G0,VK9OIJKN]+f#g11H@)a3(059/U13PAO6-(V7:8B-:^L_NAT-K&ZaNWHJ
:a]VB\bC<P9>+5ED6_WE.g4FR@-YSUSLECWaW4aX-I]-4GRG+B8H\SZ6c7XLc3bI
.2>U.bCX?.U5@X;TD3BE>S(SQDA>I9;1?AJDDI;IS7&@/=<^66^EaC?9?SIcS\XN
d._)A_H<9cI(?)GeE6/QJ(Y.BD(H6f6d>U=B8JRLBf@2UCf\f6JPKFWF;=BEg39Z
CDC&A@7?U>eKB3Y25/;\dTS1+_W1YU+7E&QC=#2+YdW53@T6FY4g:2.Y2e+LXd+O
g#6RQ&A&UE\N)KDVaDU9S1W4ZC+]N1\FMbXQ;6HNTCZ6FE3bga(HA)@OI:[ARP#G
+/I45HGHY[L=C5D)Ab=^6M-2.B+\ec0/NS;(_LU/7FcJA0/c;<HZ=d_;C?/=e)[D
EY030DQF9:Q,QR]MI9c2\FQ7R8Ne#_Z3KZIJ/CMeEF8Ea^F&,D2+fHW6M)dXT=Ff
\Q[Y&ILEU5B/c?\LZ\4UIN>._ZXM,6ffQag5SJ]eg>JH-K9FZ()OTE.0G[g#Q<&g
f0\\B697J0^&A)VM3A#Ec3[7_7B1L+b\4),d+eZ&7cB304D=bZFR]BI#5+d_2c&0
:3\g4I,;,@:51[#YQNe(0\A63(X@8Z+fTFYa2@c0S:0M5WS9)K+VUZ2NX>:LC#+4
ZH0&)YE>+3Ua9UI571YXcdM;DRQTG;(0T::[Q5@<PBc^@:5UO&=5PX8gI(9?Y5Y#
/0@+2cKEA>(#\?R2Y1)2aONYXXWI<>e(Xa=bYdG,QU\e><N]VDafHgW:XZ7MH#2&
/56^AOD:7SG<?EfLV;=S2:0<GcV;FJLY6Ga5)_16((&>J-9NGRTB+V3AF:?>EcBC
[&@2]/G9R1[<\90MPZO5Wb_:7E(I>W7@:5_4^/]aD#,1>;)eWQT0VI?I@.@Y/,M<
Qe7bMcdAE(MV&?Q1628T;^XOUeEZC3UDFG_C]S\(M&N-^[=\#2Gab_NIX0BgF_\#
B)FbA]Ue:).:Pea&+<5NX/RKb<42M?2&a^]cP[@?:;_Zf\RI\d:>G^&R/\dV1>FP
Yc\UK:8@#\fY4Q9MRPZf_Z(?ILD(E4E+dJ4g9b48b7aJ/]@4a>PE-g(06^eIP>&&
.aNOJOP,?=VOG6^_C9;@82(;1=.MO\He(RgU=^;]:&WC6?;59M(GY\C6H9@.af;2
0fb#19SO.7V9QRI3]cC<^ZVd6PTC]/)aC,A@.\MNICKfJ83GQ2gU,ZF,<2<c0aLN
/?TP5B,CC)#1]Y<OJ68UT<.];LUMYBAe5+d4==7X>U\Y_3)5SfN(?cgg_XYWK2d\
<c^W4265/,M<95UCF7N3?K/I@=eX+b8R]Ib0Hef:.a8L2>ZfXQ/d6#g6FEI.RRZS
I-6&1bT;>[&&F9SaD@-^_)OHC59@U49Q;J_/PB<&ACVC<c9-=(DBCcR:>=eg9g>,
7KGQ_95-W[aJD)[c1COYR/I]O=eI,.gQ4A7Z86?=9OUaV4EP&CF[f[0IU]QcLB?B
:B=0^Q_2O/\W8[G:0,PeI88U5[65KE81b=Z<]^J.7d&a&CGX;@_UDP,\a8#AGEB/
.^HI=8@Cgc#@T[?bI.;)@<A=3]@-V-MdCRK#C3#-^^O/E]UKV;bI:T=LfcE<,3#V
_#Y-.bCYe0YfE<SUda]?(eaP4OCC0?aB8U(;E@LRI=[<;R)L^C<(7-ZJQQ0^1FHE
6U=I/aM#O0>)^5LUP#KK[D07g@)TCT^;YFMdOX5I[9T\3NJO5M]:D#gHZb<=1aGc
5\,#)\>g<bL38Ng-f3O]=W>4?b(Z+]WA5)N:K]:]+7>&//MXb)]aRBEaEH)X:ZG;
0Dd\PJf0IC/@Xa1VQa>;4_.))V70f?J5\ZNXW\IQ4-^2;=B7.+K[CJY#c+V_aUMM
7LX;70X:#;95HXA>T(9/=OS&BcR<6U5;8/29N+V&<dKLY7Q+,:^Md>B&0-&K+,=)
?L><<A&NZFf4g[N4H#-78D,<3S-]C6/-M]^@.N>&PX:_NO2TEb;a&L,0L)=#Nf+0
Ig@]=H:b0VdAd:IaP2#Jg/GP?3UeN^<:P)2I7H(<_CZ@0:)R.@=TEbT[>g;/5@Z]
0W9^=B,>&0@fCI:8V0Gb.FNWP8ecHE\;]Y3\<(UXU4ATfZ<N&2+Z((VXYQSJ65+,
TdY#<O]LG)gHUD01-QK<O1Y+UJ[8Ug3<>Ff9TX<0RCR)/ae/?d17&,0=Q@(1::=B
OJ,:c\:f:;J=./[P7J9MJb(&IbdAQc4E_U90.f:T9gV^\DNUgIJK@Ga)SE3R]Gc5
=.V>\]Q,B<#FP;Y=)U/[Kf1>0T?Oa_OLAMfbD#X3:T4@I9O,Kd94:H/AUM]XdfKc
Md:;Ja7X>^L8cM>\8#@749cYdVR&RY&1[aBVR+O=Vf.B47#4?X\F9P?7,>egA^VJ
WWYHPNaZfLP,A7R-<Ka<;01.CQMT\66bK^86_IM[8VTCHVMZY/4_.LU4JBc/J:d/
?]&0TOFPYM=_2:Uc9I,)e0XaD^BHA@g,R\SSBMP/Z<d5;ZLG.84K54[G<a;_\N^7
2)^KaJ(fZ5f?BFI1OYVg8IQ.,aM;F/><CU>BLGM&c^G0g[]#QVK3N&&>WBc]a).]
T\#bAaHDT5TI?6?T9ADKH/6cE-K2_J9faC-9=Nc@HZ1)5G6TO,SON=CZNGR<CUD^
MY8(Y+bJ?X8[9.f)OW:Da-I)3WNF73DA-?\^^a-73dKRCPU,#5^A4JLB:^2>Y5E0
PPgKK1L=c?I+=QB9f;(:K)?@2]+ZCGP2BgW_b/CX\M^BdU1,gYIV9L+f8dH?F8\:
XNgV6A,X@A&OBNBLQC7;F[0(cA&O&40@@B7IA0K3IYSKKc<BM.=,#B5L=4]c^TN#
\dR&)LZ4#dOP+f-^5?>ASDN:>#Lf5(Z_:,6:E5;@L-Q8D)&@\Y<N:D6TaC:60)Z0
GAG<,LgKee0OU[[WJ#DZ[L[?3TbAFFP(92Z1]7aOVNB_UI2^N^Y&P\:3N/LLSc++
A].)I/@LS=ZH960&#+TJGB=KY=<(cWQPR3-=B8NH+R@P7W:;+?,0DA6<dgI73&@?
]fKO:AO<+GOO-R&1OD.(\@E^?8]LE]I<-/2:[=348K9K-8c6@\bOZWeL?&\Fc-<T
?7OTOX7.ZRT_?@]L;Q[5P@S6MH3.G(eW;J+8@)D1I>ZJ5I+:_B1=6=D?,:O3;988
:93GFX(8(659B(GO\6<c=g)Z]GBCRga(<&<;X>P7<EP6)I_\35EUQR,Ef(83e&08
X7Y835OgZed)S>YO)+S^dO;]M3(:8T7A67U1XUSaXf9<<BLS0A]8&L35,IL^_-e(
G#<L[N]b/6,H5^B#.X^a=b.g.Of5L-F;0d)L\ZQcI9X3bUbaN--<@T--6O)80gc+
d#OHDSA[(NBdaS)P0gScTMAR/&37cLI>-JaTB3X)3A3@PbDE3D.T-SU8fL?7QOHO
aU#[I0A=,^IVU&GW.RdG[CU4>#6#036UWc(aD3+);XSIQ;ER,g^9Xg@f4E:;:U<W
,RW93/EX-K[)7WM4bK^8-&Q^bSUT7gR[18.\U3P_f&WH\S;+AZD_9HG\M1Dc\Z\<
aYKVfTf/UHB2SYFf316gN86)).egW9264E<OG5-[gXPB^;gBbA3AZQNd>V9\.X#@
MdBgH95ZY4JXDRI[_3ABN,90NP-^.^a0ZcJ&T;5da]O9&PHD@<=@-2=,a2_T/RB/
^AfU17K(^OG0[#>#051C_7cc:7Ie]W-Y5@f3U^6M;8IRR3_DL1gTDb>4=B[LA<^g
&>[Fb,;PC9NJN_D4;:N?-XGg))24\)B(.PFf0RP8=1NOY,.5B[MZW-3&3C[1,;9&
AI&Dg318/C&>1GWB0>;E1O.NL>#TU&-a]Z)^JL(Je]49:A>@82g9IK+(MY,,50-1
<eDB&8MMN<3Q.9_IEf,?1Ke2U,8IT:81]5DR6.GfAR9.Z9NS4U/J)9M:9V0#^,dO
_E53BDIeJSYRbJ;J#)dJY[fXC/TaG\]f\M./6a4MT/?U#6G]_fED<f)42[cVK@Q2
-J0<MH0FaW]fPQ6[UBC=E@d\cM0-WLbac?(#WaL/BK;U-f[Z#(TLDN<f4K=/MY>]
bW/MAV88S8M#.KWOINggKS/79)3E@9.OS+PNaCgD:[=;R5HJ804D#P#RX;3dFaS4
^U_NT@XMCZa9BaT#]2HJE6L0BW&4HDX(1D4DGEI/G_gD.]dcX>[Pb4--[72]f1<b
>b;2_06Q89BRJT72+4(L\<2Q3U96E2IVRE?7DP>GbaP8O4+MaSK&fKTe+44cgbL>
eRQfH/-X?@ORFd.;c#3UGMDR,c]6P34SF]I)-RG_&Gb--YHM^,8@M#G5+3V)G9DI
]370N9TD/=:V,93S9@QB@9;LF:Jg;ARaGEA6#G65GDF:QJZ#bY_EUM,Lb>]HSK6)
,RR_/a[7HKbG+6=(KM<3FN=J6##WFHB\Y)Q;EVZf=DZ+&0ZV<I#?SKGVINbKa>f4
@13WIK<[7PA,?EX4Da<\B,b_a([&1IJfIcS,BZIQ.G9L]3NV_.YOU6Z;_6e2.bb=
,e3L9e>M>2eW[Xd)R)=QEda^31>g/82c:)/SSP-W;-9N?^^^L2ABd?K<H3MgQ9E?
A\[INJC1fbPb3H7?0JHG((=J^+.\K]TYRg&ae.g.3O=8L,]BW4gc;Z?[TQ:f#\;Y
:Q6Wd=KNDOH3b:C:8Y[,3./N:?]>,?O,7=)GgX1_&=;CR]#>#cO6=P-f@TX,eXIS
P[#W_;VTK-=E1Od8;DMFd?FD;-Ra^5P<1]/P)c[AGV=5#[ICH<#7T\5I^R=GMNC.
E@2CDXVM\0SG86IWLcD1@GNGQJ]LRc<VNbHP<Tf/CV2=<He@>A&RUf+CIRPO:a.U
)L55>KJ1g=b2EAVf;?4[F[UX2gQ87ZNPa&@B,><W1)&PH_@E,OOV\-1C+D/G2_;G
Q,1IMW9L,O=?ATaZZ>PAJB4QK,TH1:Y1g(-:6GRO-BWVe5e9<J_QHD5O^JJP-<7I
0e<UbX[4[,-8E<8>7):PM,0EINS7KF9Ob)M8S7M#2HG7Zg5X#dRL<1a>65+QO\J&
]+T4<TJ0I>W\,+gM4<-E@S?4fP1?VagB2O:<V8#F_7&[<VL:P2cfM6,-P=F^(D[B
O&]dYR<UgE_B49\.Z_,\U8[JIK>;F(^^ORc^F1DNH?\?DfbL02DU9Wg.0g6Se2/=
G_+OYRCAa92Oc#OC43(-3VLcNTUIL&:I8P0:3MQNe<_R^=W+R+54(1B^D>bW]XHT
b<g12:]I.K1_E^?50g55_cG&DW(N(dG3SF+/#c58ZR5[edV=]QA3d5HWSGK#e\\F
7NK.94W@[8EDg8:N(_<,R[DA=GDU-d6DIIS.SIN59=gA58VR@GDUOC3ID,GW6CN8
B#d17DbS5GRDG7edF+dOE52bT)&)26LD>W\P)W=T(2c\8;Cb5CT_I9JT6/1G.CfB
J<WA@TOeT22E/e];@ZeLRT<L7?SZ^R&C,VG\e,FXR7Fe,])eW;Y2DXB[Me5dUO(7
<,GX?;CT[DR3dZ0TfSWC#NE5@1,N10>?OS5.=:HS]KSb_1_(1>W\\_9BD1N^:5g,
UAfVMdDb]aR]J>8UTc=OLPFX/Yf5d9U5fBVeG_WEJGd3)@/8E&0WDNXc>MHbTDG/
:[7VOW,[3SW01cc9](Y>c_\;7V9TD19]S=^5cJ17&A>a5,7,Q3aaBM_Wf(<CaIdS
RCGcF_g3g(]E5#Bd0Q(/AgI2K6RNZ@C1V9R?BJFTLRe/VV7+:P/D@0:UP.Z&UMSS
6/f9^6TK.2XcO)1UE&+FX)e-F-<.F5fcWA<,ISJ5+H4cSA^1\8g3/G3\=MJ.1ER#
@V+T2)F-e^=^]VA;IC1d:+OXIf1FDDRG=X#X^THeRedEAU#.6SWCR<8.P2YED@Ba
W3-^YK-MQR1SH8CXI.Q5bNJ@[WI498I2@#L(bNJ[:#<)FbN,,&5@9WPA+:ZZ]-,4
FaU>5RVJb.&e4)NF66H](9RC\TE,662O@7N8>@P)?U/YVF4)dF/^GEA5H,AA>S&:
6Xc,ObEYS8(+./ccM\#J-D].@[VXPJ7YPeI^[_NbELH6X4.[H)H;QUcC1>Xc;_]+
4SMMU+[A?5F9ES.QRRa&S>N&,TB=@;?I>CF94]@)YHLCgPZ#CZ+WcKZNR1/._>H+
-4BG\K)9P\_S&(SOc/@Q^06\bPbWC_22aJI4.,f6_D_/3aIXKHNYeK<g/NE\W;F_
FcFOP5B5R1QG+>&L)DWeO_ZP36S@RV:9CfE[Q\5(Z(IHDH3]40@a7^6M;CJ8+8>/
939C&P;E6<[..^2gO&I#?Z=/cW]B8-e\WHVZ.ITSBdcg3\gD0FcU;IGRS1@dV15<
#gAQ<fF7C#AL]C,bQ^VgE<1;M[55#C0S-e8J(;Ud,\/W9_O4^=7J645GLU(9^I,S
H1=^>[?edDOSM&U-6=;N9eR(@8-F@P6Y2K:L4[DdWeW<@Q>=Tb)OKSQ2JaX]4/BX
#a8<SC-HfaP4J\OB8PC.5>>QE-1>;X]G(1/><9,;0YaO1G4AY.0ADS8bJgJ3b/e#
LQ)XBNJV;]@H&J15&6)fWIM9/4Q:LC,35CCYQ&+K3\bPK@\dV5.ODWCaA>JgO_5;
Q9)G.V0&9(MRQ-G2SO_31V\L59e]V5,)D>4bCO:&-++U-:^6;dG1,?UF;[#WdR]:
UJ-[<#.WJTcJ[J5L&2_[:S@8,L#9Fg09.cNP86QT]&R8\c(AP?6Y7>H?PfQDS#-I
#I[.MOb-+#BAB@Zc>d.@AC<_)ENW72?M-aL49]HV<L5@4BKU(TXMac.^(a#aFV_7
c=b39(XM#NeHC;/+=Z@P.G/eLQ61UN4f<&FaY.1>,CgJP>LdUV;gXbE7SE6;Z?L8
J:cDO3@^7UK(V]ZU>PS>XM<(O0PP[X1_?0bWe5;^feT7U;5J\gb:.U)WD56@d2>(
BK\K#TCIUATS1GN.RLeNa0^f5dQb2?-FP(FWfZ(=&O#6L74N#W>@bTbDGQ]?0F__
SQ0;N0M=WY4FGd:(7c;#78=G2NZ1c??ED<T1L/TbUd=e=g\L1QRODX5K@YM8R/e7
f8L4L[+=66eeWW9C>1c@]CD8PL<eM;+)T,M+5@L5YOUTZ(F@+O=T?Cdg/b@,CBH?
4[=J7+<S=UN0d+]IDGI@52NK\Y)V5F7J)ZHaGK(->J6;P]B]+J;^EL1)#96W_WD?
L0-]B/[#Od/;g>I0QAaKgEAT-_D/5?6bGO9L0:I]C@dR^]DAf[7AN>GP[X7A_4.?
_UeLVFcbMJ+W@1X,AbZ;R1.&\g#,Q(M@EGf16U_ZX>ITJ-8HH\/7AW1e(\#@84&)
:\DC?:4dVF>O,T;NDUOeYR4\TJP3=6K8W]ZZ;C#4=0RG_CK_&acI>R#9E5OBDd--
8&[aD^9dL]#6WL)W0Z@M/_NH/QPI\aNECeN14.B?^+bTg\:f&O.7@fQU69baC\PH
03>cW_(ZdJ14/IV^G]+.78].2M^\DV]830)ZF3bRUTS-+N=<H4?;#=&#;/?O2STU
--#U023.38cZWACO30K_]P<a)JTELX+(>B73fMe;c&SVPB?HB+N2GIeV_\cZHaSY
K735U22I^4-88&J[AH-Zef]5fR[?Gg\-#-D/VNRV>2_dcXC)IZ:5ZKFg[7P;\^8O
eB4/>3:/>IB-0/fdYdC_TgNS86@J9=XJ9Vg+U;7#7O?Y:73U6D6Ga4#V:>Id041Q
5P(9T53DOdQ3aD9Eaf]>?CYF_XYb]<L(-f)A&ZSN.?973<A4<HY,9OX]CPLO)_(f
,O&=7dXcg5b\3Qb)?A\gGP5<e<Y0K2YBd#(Jf4K[]I^D+eJ/8>-9P2YO55.#b)-J
X9NMBILY=eeU4J\:g)57H#3E\XNHLNVeT5.K8J#f@?+3DbYE7GZ-f)AQ92QL\[?C
6Sd.HM_2F#>BTA^BT4V4-&bB9_TC)d0CZFQ)&/@1A]dfZ)R?GgGPK_f]C[-U3^[.
8\,LOZI]XQW9R581WYYYL1WJ+UZYfMFKF6)cc5X2d4N81W:EGX/QF?BH+=N#NU9D
cT[9I83G^^^BVI\ZAX0FNZfP&eNdA?]^FA-.E[ZdD3?HBA;.#TGPa1RU9P2>=)GB
0[?3,2/L9dBMBafFd38G]-,c.^D+0#0bW;;]=d,WFYd+^GQbbcC)]9d>EQOHCBKB
)Xe(eD[(Y:QDELYLW(8c?@(HO2QU-A.N#),/;4,&E.U&Af^:<ZdJcQ4K^ZF]C2=\
Bc>E@E7]g,U]^S9&/<R)d.c/N-[b:V@+Pf?UXL2.ZI2O=+16WR^DX[3#:/4.KCN[
R;&VIUGBLXJf3e#09Z)fP?c,\/JOA:);A?-R,9:b-e[gXg(YIf47c6fOSS6,Q-8X
A#g5B>fGG#N-]^XX4K+:)8Q_<#I#^MB8b8bUX07JV7QV\E7]L81,QGgcK:<7>S_Z
JC1_c+6f?FW(GPK(c#1#1TTP#J]?cA^g=dIc]CUM-1QW-A91P=@NI+Ie\T0c(:MZ
CfH&?>CO7-;H[KGZ28[1BEdS_6]bHa3=aJ[\AJ)NJ71\/&W&OI<1\73,+@TO;(1B
Q7NM&)66+N7#?OA(HX4V@fO:773a&BIe#+e:<fFXH2E4]4#Sf?<L5142+M.L:g7_
8J[KS.-^KFZ;@&?L&g0d\/2HVc@(TX<9CTNRO9g@W;:&,d#-F(1]:aT<XN-0U#EL
J2_3Vg8+0BQLCJPI<V&&@VDJ>1ULFe0Ybd)aLP<2Ab)-FZB=4-e=GZ?;,U8eJe\e
J]#P7WfMCg5JS9@+H=LZJbXaG.e5UU/Z95;D5cOR(_Y[UY+AFG[LQEV4ZD82NI:Z
K>Vb5g754#19TRE&8=F.5[U8JH8<ReM[FGUP6BI0Ud?R\5]7C1N+MWXdB3EEL)R?
H,UOC:=QODQM=&2&[\b2_LQ3Z#Le(F6;-U_T:#8KX3J(B&00V.8BKIgOPPeF/96;
GE,UH6\V>90@O_8KJJ\8gR-Z/,(WSgJg9G+&GeJaBI^301O<AW:/Je>=S+Q2\LC)
c^aT&)&NHFYNE&JD;+V=X+5RTW&F<40J]8)_E^5[5L\G@@aAQTDUTgP):Wc+[WGP
@;0LA]@D0a6:B#1bSUB]Q0=.[?#4.)(CfDG5TK+4SL;S/#4ANcH<Oed9=BOLcO:g
&7B?F@M&:+QO\bY[S\U.F)VS,Ye:e^^XD1Sf6#9@BCf<5\Z(;HPWdAYg-=,^7a)F
7C/&7[NZ3Y+C)O0+eK8Q9g)9_eJCKW9:8]2XZ?]NWeD\#5eMMPF2W>Ub,B,\+YdJ
(0/,?:7SKMBJB9dJQDNL_-?QE\ZA/b-Db\MAD?fd26U]\.N#H?f2f#+/-<c+O?PZ
a1L3)6?1decZgO,aT=[:/-6.,-Q7S=&)MD+.74eSNB\[P&_)4]b>2SfLAL[G-JQA
BKVdC1)(dW]1eGZCNA]3@F?]N7H4Y:#PT@[DHB&#R+#bf2?F?bPI26bEKDR98TSa
\/1H1Ae]OO[7^EH]W_EOVFK&)Ff+c\eK8PQCH(#gc:^?E+S<3KP8R>;b@Ka5I\IG
N:O:(8JgE>ZBg_:9fUO7+gJ_7[#XRaY,FNL#:O#/I@DHNb#/8J<@=P8fNN97aPTC
.b9e&FC<]dgV^a[./36>_XZY54J<NC4,d\Yf@_d5Q#DeNTH[a=/3W)-5Y^f,:HA2
\Y<7P8P^;QL2T+0>DXf+A3BMYK9@D:aXH0>J_C,FA7A&;2JB.:L=C+<f\82.WNK0
0,924=N1++&CX>d<93=#]NdB(QcO_+PSRd2/Q)QQc9fI?/a@cTe+I?;#6JdcM\D;
2?=.DX)_Gb^aaU)X5^55b:V[MgGS>6VWOg+646[ACR@SCV<d5]<LHRDG>6Kg7@CS
Kbc),6,CSeG]5NOKJBA+2CO2g@@d+[,,J5HO\,-12\/Gg9A4+-;NT7R1Z+/+A,dH
26Q^A99\CfPG.U:UO^cV[Q#LgeEeHcfe]gXD9@_aB?OL7JgA(VBZ7OFWgRV/CB=[
R;&R1CU0:O_4O>DB/<TKeS<X1RBSCOLeA4Ofac<f@_S42+<B^9/3O>T(.,dZZf:9
1<HAX9QOU)78<K_fJ90E-+FO[E#^EU3T2C76ZaOX@2W#&a^M_STB,^5IO827YR+8
#TdeUY)7V:0,Z8WNaQ6ZdJ-?]BK=-g)?V&D2^VSad>0Z,#?USPMO.Q=S_TfHaeGb
EZ)2VDQ;_3,MJN]?D76<ECKe0]P:)aVgK-#-;?Ieb&+6>;cg;MK9Y:e.)ed,^a]6
KC\S02-4,(RDY-K^;3^Te;67@9/Kg(+PAGfUH8L\9+Bg-#)Z]4/DJ<bWU>5cF\RH
Y6S_B;[Q96)X\g+9@.X6YYbE-+EJA=L7@bNZ(=(#Ee+G&+e)MD-1PR:PS0\;5a=W
,\bRRK=X?O44GLO2.UH9eOTYI1;O=O-IM\6BAKgWMH6:9E?;?>Z-a]\B;ZP-4bf>
f[c;:ZNOX07O)<gc(KVI/cM#LU7&00G<=f(f8[R@aeSH(Qf,OM@2O2OEJ.Z0;A6?
1_]bd\B#XMEd4g&S.+AK##6C=]B5M<b6,.Vg/Lf?=3XdPSBUL6UG+#A9YFE:T]DD
64\/=2,3WE?3TP,ZDCHfL-EZA<Q6_UR?(V\X/?#XE[H=(7)X=&A<41].,>BaHZUY
R2J,S^3=6b\+/63T\3:bN\,A^Z8TKg[^ac5GDd4&J]#J1LC[cMN>&MWCR3FD[T=O
(6T4+Y3#_?bd,#?U+[RS;@bB6cHF9R0.VJ@\HP(HdbFDV@4ZcJF5BEO2E1ee7JN+
0_1+1=We0f8EL##9RBNOX[/URVWRLGQIV(XLZb#Kc))(5PU6NVVJ?X&B[Bf[Y=.W
+>QaT/;0CeA)TPPJJ+Q)E2=,\IA0b8C\O_K]28:3eV8e3475:_;]Tbf\13I7WCIK
\cQC=PeT_BHMD;f,>>G9\5.:FVTO9Q/eD(V+=RaH@P&.[W6&C.&TS/X_@),;.^[g
Ye,A.WDZ?Ga[IgSa:X3JAR(Bf+Q<?)OgMKO+V.P>DRE\]\[L&LC^ebPE3WL9MZ>>
ZY:GEfbZ[_#ACLF7WRAR(OW;VBEJ=HU:RSUbQUJ?a6YCQS5@GFDH[PPP/a1dLfHQ
6)L8H-?QNJWZ)PdM?6/GX&(/1\(WSZOOW.PUOH;4Y7UF=:,HMAPW+&JKWZdg7=f\
:3_5\?:_C,M2OQB1>/)dH\2AA>2YT_b8(W(P@B\@98E:0^@?XQ.-[,=V__>LDQUC
T,9]AYD;JV0Z.D1O//e\^S=BK<O4@C2B&2OCIWNQaLU7:AR0ZI8_F>g=C9L1b@>U
[J9S8BWa4IAE>5O.74XM.:Hfe;05?:/V?&V\5OL/4\(DFdGCCW#5,/^3CI:F#Ud#
BM/F5[d=CT2;IB;@PV?FN_3:>_5a38Kb?K)[Q4QH97.Vgd&E/IeB[dMe@@K<7NBg
6W#C7g:3E8\fZ8Md2\XUdD\1@+7]M;P#,FeLfe]7FUbO,>_LDN-GfDNSdU\A4Y;H
)^<@L50Z3)OM_CS7_71,ecK]D.GY#f/@4UfZTMROQ;9QD/4K=<QP8=U?.R.IWaY_
/I&-:J(K3\c+\.a&RS,R.1S&[TY+9\=CA50JIDY0&(IAXY(A(FDbR.<7]]KE/S4X
U(150L)X=B0f@aG.GI/LO/T+SOBF4):H6AJZHF9fY^G@55K?F.O?4CT1:]S240D8
[<3(KGR9C[4RDD0H)a8f,;GF9+[)9YPXL-N9(G_QMRL^(Q-WEQ8H9U.,#Q50_aS7
4aB\-1QQJC3U>dVPGG1c0PS_cA9KT&DTI6-L1I9]NSK\1KL(M@V<O+@e7KNM@9[A
4gbSV6_-U2T:[&UN4.]->U?E7^PG@>V?/d-#+V&T23^KJ3U-6<AC73NQceH.C58B
[#@.CV2CXZPGe@(g06:a7c=gXE<OBZP#M/N=.W&^cD2#g\C.\K[8HK+8(_4Y[)\[
BI=WFOI-c1T47V3.XEYJ:6I(B,CM5<I@WE(Bg/f>W;f\[;GT1^dEM&ROV;,RgaT[
832((>9?d,dH&?;415@cNeeB,cS.9Q=7f0##_1,7<_4fV91B;8e:bRBJ1R?6fY]?
R^4?X0Mg-53c;L7B\eN#J2\[;]J&,C]R_5=_OAQ)C3&T\gW\Ud,))MLU4a2^g#5X
Z+\/(gMdMP+e2NA(5BW^;1X\cVOK##ZQBI?4[YX3Te3a9OS^eX64G_\A6Q9c,2<\
ZTX(GaPeA6Jd(@MZABY,YQ?OR=1I;GDWEUFM8P9cE0-Q)9H4.V+F\Hf8cOK7A^S1
Db5W-G\O<HN#O:#bY:&<F.XMY1LLD0V86WfYA:]P?JN0K2490VA)U,EJ;2<WM6Z=
?J\Y4XZe(\9N:3<Z<9G=->3fU8Jd7_Je?TB#S#?\3-a5<W,fCM[>?L,_dB/N@e59
UG6H@\966eIS[eH,d#Q4Y8GLN.TbP:C_c]fM?eAe<H:G..O3SV0Y<:MgYcH[G4#6
[+5R/(?&9E#[_U/OSCB9._?fBJ9G=Z^Dd8BK9eecBg/A2J902Q[>22V,.:8;IJNd
YRGIc>d<QYYNW\Y/8F7;^A=N2D++O_J.+Z>Q5\EUb;P)K.a\5.6IK7(g@T2(3=6a
\(1aaXDE^e]#0dP:(_=5XP<-TGEE^2NV9b(JCTS_\X5-bFTg66F8XK_>R2)I@[7R
^ZAW@YOTddJ+:I(](c&GN34+\@?OYJO_La[LH95bR-6#H5&.D>L;;=7MG9eOb\62
R?3X59QD,))^E#Cg(N0eI04J9E-P3@d^Kg5O0)&41,KA<0U,,2.W3CP.SNf2(YQ@
\;;F7f><:ZW\g=G?2/94bBTMX7E+bc9YD9A+K=12#XZCMaVf6W1X0?4fd<E^03UD
[.AU;-F7UMLP7XJZ-W&Md]06AbbP6:bQ&\HNXI.@d@f[e^X:2S_XA>A-E_=cK[24
^],a+Q;,BG6-+@ON4?0]S1F=bL2^L&KUA>6AdQKfU>gCc(8H0MQ_;M6e(2a]\0^S
IT>P3A)6X-Z/P8[CG2.Pd(1a46]eC2K)=V_^[0K_R#\IBZ9V+=@]7[?QHY\N\UR-
3^,JbZHGf3V>0=_FJ2fKa1MYG&XOd_H+R5;\)(\-,@WVWdf6_1Oc[<E@;L2GE03&
f\9Zc2++6NCD26[1:KQc3fOZK5C&><eT8<#RV>g?-c37Xd>ISbbfgZ79AX(TI5Q6
Id(Ac_R7L>6)3g;CJfZM6-O#;S?+GSX-RPJ]CDY,V):e72.f4c,?e1Ea[cf]>efY
Sb8AQ<,)PW&8_bA?K:K,M:KWQL+:56G6:aNATW^1(^&F&S]QVD7W3K#?V1b+_L_T
EPLBXT+^@W_U;D8K=OOS^UJ9UMB)TE;5^Ca-FVL[Td,#(AR53O[W.[c8]eGV+80B
SW#T/(Y;]G##VOF//O++SH09099A\,a5^WM)#T;PEd4XN_-^-/918(?UUW0g5M>(
KXP2@I(8Ff6KC7)[ONf<?+UcJYM2^DW+g;?<HYAb/CQL?GA^1@dEAVQJa5-P<TQ8
/2NM3D-@#^#?R^5^VHH;<6?2XH?&O@7(LAC?IYV#RM3Z8QE)D3QIE4DLf[d<C7^a
9S:3RcRBKMEDAXK_cS9JFR14[#?)G+1&1.HGZb3eg5cWF1ea&fe8N&T@JeT0,YLY
OA/\QAJS2R[+A/T:e0Z93)_0)@D/KaZ=,&#_,+AONN>^e991?SPGe[L&6KH6c3(K
1(]FPR:6APf,gD-_QS4O5g7MDF[4He)_POfB2(?JUVNRFce;I9WeBeM<(H-HbI\0
Fc46RU1>@LC[&e,BegCJFX2I=DWKR@+RV-f\]L1Bcc7Y</>9K^2OZb07_C,;G<\\
f3MO_9#aeDfBIK6P0N_]W@V8/YFO2=NWa4<I?4@:VEA/H:e-X3KKVIM<7/Af7O^f
UH?Q:E13B,EJ#^)Z8Y36#+4F5@^]]cS7#B,H1=abg]V(1>\^2#+1@S)Jg::S14[a
9V@JO=.;C<MMdF9M9A=J/_]>JETL#(#N-<J3DLM.Ye]S[d>VX<2[[[a(G,-.:]\>
>D:eVJ+Y,1;UW+,5@I6-@V28H2FA6=QK1]G#.ZD)bMS3OPTXM3<5>)V]U0,[UCIU
>V7(^Q?@#IAC.).>T@7H)1EaMHE/SJ(#DTR@3@[Hd-V<Wa\UBKU+L(_@#F@e38G8
dD4SNbZTI(N5]e.L_DPaIeDZ/E?e;Fd:?]T2QC:J>T&A7=S1L==O-@PeDEQcKeg<
4eQUEbZIUH9@:/9;CDCSKAOWFcJI9<S<;&4X(3:=0T1HY>Ag,9T@cH2YUFa\S20g
Hg+B?ZE.P=PHPC.g@b3(gU@60X[>98-O=OU/&b?LAASR;VR[(c=@Zb\EJJW8WYH0
]BgMg;BZOL16MTIZ\J7NegCZZ(6S^5OfN#NW=0=)?7=(#6K9BXJNC2U,DcE9Rg<5
&(-MJd&+_d6(CFL>BgUI2/)g8A.\IJ3],/].+Y@@g5O,d+a7ZbG[:.cL1c7CNMW>
_C-#.6F[@(8bb.RWC_4IcYH,9Q=>gB,Zg<5Dad/9^M.@Nb@fSW.bCM#UI2&aHXOF
FGVJJ>?A(C]L+(c/[MI=\-+\+=(()+3^3-AY3&KbZRBG)5AT<G^=H\JQY&Z1I(_I
@):=R+UcN&3-JY+QS5bJ#.)?H.QM9H@KH,\:]G9eFbBZ2/,>+?]8@PXB7dgU0aWf
?UG&RVYG\@7LYg.GIW(UM0@]KYQf)b8,OFI[@^fZJJRW[dKUgKOHPa;YDX.\f,S5
IJ4(?+7b:XJE2/<BRF?2I;OA-^/:H#b5U/G2/@M@#c9CfB>ZDB/5ZEKDPJ3GFd4b
aE?T\^3cf8f#6Bd2gc0;DBc_18dEQ\B@Hd.I/AYZ,BdS?\=TgGbBa(Eg=.DWSG<X
6eZ3VIe?P.gfV,SJTOA[ecCX.D&R,:dCKacR1#(IX6&G>T4-L>\RVLTG?O)^&VGR
3d.+JUC1c>10PD&@bKNg7:P)\/]FSNY(YPfgVMZ<-g\g.g0IeGG&[:SV,IQBYNOa
;N]?7(Z0LfZ^@#4ae/2^[8M85.7bZ(E;OOd.L-R]GD3D1QbXFD=Z<?CV8?^dQ,E.
U?d1>\cY0eecMB)aU.:Q&_H+G?K>8NFO-;KSQ3/@VRBH4EM9(;1D2^O>9X.8^9g;
W2>:7;2S3>5YG_JcIM)F^@M\e@:Z/MFO0E;&)R\D\CT,&[MebcU_8YE&g9,B8D9)
FUF\1QOYJFKH6f#VGR;4Fg=+.Q6WcdQgN2g]V57ML]6\(dP3J2JT@LaZ1(NZ?@I+
\]CTB+)PL89:\+L([1PdV(/7e9AA15>=O?]/fT^SC5HBc]a1NOR9=+]>R(>e-^K/
X4H.b^f2O[Od.CXV?^,>#N=4-e>-<ZD4^:>=M-/^SLU)V+EK+f?HK6=<]H7F(FH>
VR4&J/\@g,SaK/2;f3U18?Q8G1<R&YMcDTL4KAI<&bF6aS>G.&@YSG.V?3KQ<:HY
52T#ZgW-4:dTJ0:9?I;NO\J?@CV(IXgG0=U1BZH8a[??.NbZ81(#6c=9(6<559]d
](,H_V#Y3K/5C:4@_UIV+,)Ac(KbE?HV#]?2f27+RQcc+?:bGSGE@+U)Sd>Z&0\7
dIO=A>=1Qdb-[J#G]OdcA-Y@(0JKY_#0+(D^(5[0Q7WK4F1T?KNe7dLBJ4.I5L0Y
_I]CS2[OaaQL>f67I3S#1B?#I[X</He#&Lc@Jc#/[b3D>TLH\VIBGF=FgE?c^C2S
A4R[>2U9NAEaVWTSYDe?B(e7(DCTDI>L),,X7W,ZOHfHZSKWZDgeMI4][e2W+,:2
V[@PcR-]dQ?F4H863O6Q25,KK<6aJf\dU#XBWa(RZEcTLC+_.3Zga3J<OX9:+04:
bg=ITc-]JK@?TCHbAW)5>XO7;W>6e86A.OU9UFdKP2X^W5/YJAE2)AYT+eEZf4>S
Vde6TO?TT&06YY;RXC@@7J,Y8cc+^HKe-^Vd\/Tc.??#?H:O]QLcY]G?O06X.#Oc
6@+8WV]HH]Y=2:69g=-6,gbO4YRG9fEg,g5JO7bI?-U9L=_PV\Q5:VK9@Y3F(egM
GS5[Kb&M?@V)\02;JZdF@.WBF1#aK=[e5_99;7C08;/\XB&EM.1U]dM)392(6&Sf
S6B,]U=HV,&d>a-^LQ^aX.S3e];A9dR7SF;bI#^#C=)K(5EWdT0IAd_)2)RK.GR4
;I33T)--Lf?7^9U+[A.8bGGf_DBN1<J0[(;@]7Yc5Z?,#N<>ObPDIC>+OWf[\e-P
10fC08<R9ZAY58[]UOHO7Ge=Gc&J<eP,?UFAB,Q:-+c_gX2.c87HgLHM9-FNYO_L
]43QH0LSTHeG3gd\3N_+^#?=8ZT7.[P:2RPVJVT:<^#2g:CG4\U#C[RHZWPEVd;G
Ld0dJ9RHM2&,1GPD^;T6+K.D.&Ug2UHOG,?\B,f,0-IBDLe__VU^O^FQ(d6&T,DZ
J95O_/(21N=eaf)TEc\B&@XTga+L#R@H+_U97D?QTbS89[g7S;IMd<VQ#WC[MUa;
G]PEUOT2GM63^F?b0L]A:c=O:Kgef?RgK\KZ1L6c]:S4AfR[ae;&3G9.c(I=2G>b
_JB?309EC@:C<+V5dA&+^,d;ZF2XYUWN94Xc]8-B,N8+J&BUeVU&A(L:<N\aHDbc
W,V9,?T.XCa5E\WD#;4(+^M;L:1QQf(OPC1_G;N0DE1MQFRMG>@_RR.8CHI.NGU@
C^_g:KeF?_e)C=;5O@Y<dQ;Ec@FP#]3JM\T);^CY?32+JIND_bJeTDIJDbPWRX@g
bUE?/8NeC.2R\>Mf/-.3_.&bORNWDg,,H7D/fZa0NA[AfGBH34_[d:U9E)SYZ:W+
NWJ04T36NUgfHU\=.T6,(NP+PWPT]U8eAWRN9TOCH\V,I]3S(5]8T&.aUF>TAAP@
fGeYg1&b^B&CLbcV&8]@^,B2UK2?&cKFU#HRL94+_U/5-V0S)Yb@_S/b(BMW?A+9
ePV9<1E>;K6+-A=Y.TIOdRRC22:/A6gfJ&9=E&25g=KZ92gS8/-^)_)Y\F8_3#+G
f7_cQ30DS^K8IeVBW^TUI^]UL,)bG)\dZF6;W.W9YXZTQ(REC74<?=1#CX-F-UFP
2&68T29@dAP:+eX:5ZEJ=K,Lc+R5]P40KD&K&G8HMBWVbVV)E_]?N4^SKQ]DM:Y9
8BT<+&+U,e]1/8ddaKe>T.[FH=OEC)7X2K#F(K\CbAcAMaEJV0c-:g7b@4:C@Pa[
Bc9E26[+ca<B[gDad]89WR/E1Yc0fJaA0^7YB.W;\U35_(9LT8;d2XO+:U+N0))D
dO8_Eg,,&Kf(8G]^e<M4@V24T[<EG)]_4N3/>O=?b5:/6&1?)S;2>.BLV,ESD^JE
+W\6FK+eeN7HK,#SL,YDDCRMBIZP+S7(H1cH6;;ALA=34faDJ6Q-FD39e6c^9T#Z
/RX:<TK)fb3UPMd=WV&3ND=BR/&XOK5Y6dVFS+D)W4JHW^\3ZgFg@a96I=Q@[9)X
Ig7c,=0N^&4fg<N4bcd2N\(?LC&&SZRB-9fQe[(8.^_H5H/O3cI-[:N7d>Qd)8KQ
A&SeE)+N)\[ANSDUE8S;gQ_#CQG28D2MB6.cSKfUGW)0V0V[<A,f7X2Te\@b.K1X
)g(,5;d60FgHPDO0d4]&36Z+^WN1])>[#FJX;1d1&f1KdO\R7V]G1XC;IbQX?A]c
-?ZPW(#+]#):fV)(2H55N5&a7(^H41\?>_.B^Y]YFM>..dG1S8\+>b?>\FEb4_9@
0L5>N<7_a&K>#<4B<\g56U(AIgEMXQ\_6^7G4^-#f(4#:_AC5;CcTN_4)bf_DHWB
M;.P7O/Kd:?cFY49Q?c&#44CH./]L7\9eG+BJJO5M.3F-]G/#01(B>NEIEcSPg^.
D&.+g5cXZ=aZPcXO:7IQSR.4]RUJ&ZfcB@HB6?VX1@OGY,E8ecRWR_]C/#/@M])c
/9Z4&RG@8X>348+](_SI=M0?aL.9@@B:;]E?IN_T7B4X+7)62<T_(GYe;M]LYP=a
g/PX:aZ8=M9]]a+W]5C7]/(F((E;G>^5f?<__]N6f[bd=aL#fVKZIHJ+BNML.QS>
D<SV#D.\b6@=QLW3SKW(CIY.g[5a_g(F)I+b2X3Rb+c>=[&;N/(.==cf<(,YKDR1
FBBS4X63<[[21:/(,W1DIQbBe+f/>?\WFAR#\>X:M#S8N#>0[ZQ/_LT_MZLIM3e:
egW,G:?eU,UdTO&P+I[Hd3YXP/P.01eBIT;eXRB@]WN8M_26-._IIX,:88553@(=
d+:4D<4\.Q&V1d>W1ZS:HPeX9AK?L.)/4TQTG,aIZ6(Wd[Ea<M;>,AF[dGZ88Q#R
PA?DOg.9^^Zc;=VN8eT6f0F0F^=PG0Xd@f_H:6O2#N,\J5H7UHS#2)2a@C8I?&5B
.ZBL=9YBb7?B9OSGPX16>FAI2,Bc-<N.V<V[ABNPERTQ?C<CONXE^/J/Q5-T#YFJ
CQJV5MLI3@LKM4VRI(b:-CLDEFMT#+S(0Y;_((UGeHB^W[4W^WP5<9XDHS^3<87?
V355)G^L=-:Uc8FUUJ?=ZQJH+9ABW8Q.?6_C[[a#V:MVVIL^NJ9^c-Ua9R(JKc61
S5U4[([7(6]Ca4O>bUBMU;)5-A]94050K=E+W.GXP?7XPGLNMBRfGP6K4./XXT9E
>FVPY;MP.dF;]cRc]+CXa9eZ#aU)0d76:H\LX:KN.IYL.,Ff>0)L6O+S,[B/7.2:
0eB]LZDTbbIc39YJ4g7&<Cd1I8S:b)MQ/YGe7<R3W,e8P;2J#g/KG+QBFJ#:)QIF
;<Q3QODfCC=SC3(aLcR13gU()dM\:6+MN0?JZEIAF2a,<@/bEfA]P6\):JA11BYN
R+)ORbEDG=:6+:/ITe&WEHHR?&e)<&#=_^\Xg05-;N+^c/dPWU9?[FXN=-[+CCbP
<B=6Z;/1FARK]N^V0E^YV?QXS<A[^S/C]0,P8[XL?d[bMKL1)#9=W(W^[g<d:&XQ
BICF=B3=9ObPb1a+86MS&U&Q(?aRHIR8c?LX4bfJcag6U?e-dV@,dC4?(?7IWDOF
1f3V/D8(fVNIf&1CL=+\U[&]U/)K<W_\7N@JA+(:f4&bT<:HX.5A#R@_DGFQDc@Q
=g1a1I)379M]2Q<b.V40V0BQ7YD]^=ENO(V:ZOIS>41dS#_O,^>;L?&4LNdXe^1F
f41.E+_(+2UW7,\\[]EDM]3f)TcCa=W1g[WNCS9-cc6Y_;c@71aUFT9(/M4+T8JP
@QSL<aJ?M;F>TL@]S45WC)0&0)\@Sf52&8/2[Gb+YX/V/.&_2d@,PcPB+>UAS]XS
<a78b1_U4L@ag1KZJ;[FX3HP(NLAC293T7g0+8gTf,d0C-I2RW;@YQVRV9.K-4LB
dS/?JE,-#CIAX@&[7fQT6bXD/fSD2QY17c\K?2Y8-IR)#4(&F,c;Lg+6M/H?:\KU
05KD^MVQ4beV^HeC.(Z2-d/0B?\),G;VSc&3:>aBf<e6aG&XaIN=IB-IE+(YT+]#
/N+#:K[YN/0OKE4&fa\Z#CNYB(6bCT4#17Q032K_.;K5gWWeg4-NISg7ddU9aI/U
;cF8FBcO1_eURg,g&g:VFL0N5ED5),/V>IF1-UF>dc^[[-PaD_&&^>;O8f:QZe#9
^2AMTTUD)9KeEg_df4J#;[>E_C2?8&_Y>\f<+CA11^QbW[&39+dB06QLP@Ea=J+H
CJZD7Q3K1bE<ZgJSQ>c#2+#X#)Ne:P5SH(,ND)OZ=<e_XI^-2b0BIM4AVM=_IEa2
D&SPTFSfK#>0Sf;E5?1e-S3)_4_.YX,=CbZVFEN)4PE.,RF6@]LYRJd?BYE/.XWW
d[+.<Tf-dMU>P:Ldf4^>^fOLe53UbVH;H/-7;IZ,;JdPQHNH7H,;C2CK?-eH0MY>
c3^N9d83<(9=:S1BWAXdA)=Q\1Q;D^MXVF6>dVD\e]c^9.fD14&A5,//&&5RLaTF
K2J&>=f/XWb#?6-GUgS#78M@VF^JF#AfD7^WG@5T#4]\^?N94V[@H\2;[E#+>N2a
#WNa5:I>KLY>U[:./6/d=@3-/_1.<+<.fC99RSA/)/3dBa]T#fHN,dV=J+FM^N+Y
/TM:)NYWQAGc7:cDE0\Mf^ec8da.6G3#fZLb@=1HWe/dNEI5ZA2bB&adeY70?Wbg
BH^bLbJJ#W5bI7-DSZ+?IN>K)6-1<cLW2-VKS08P=WeXd]YXMdX>AYed=9RQ\1WY
_14+@-YTJKNg(XJ9dL7,Ze&Y(F=gb\252a&,K6:+@YRGSR:d_PET=;Hc9/:[Ve2_
]Q/8[)Td)-3E[2Wa7BX)A),RESP=AKXJE:L.GDd.2e/)1>,.DMT3F=ET;6CeB3g/
aF/6e&fJXAV4bT:DBQW/.WYU&C-a6)C5.&df?CU_bV.OG>.BbYT]_d+]?(B4fV+f
Z1.Y2^HY(e)DEYa^bOeKLfgfR5f1_F7eD?P<E)IR-FO;[<+GO<?;gg\P#MYXPS@X
2.cRUcOabKd:UaH5bKDXOKS+LZX45Y\QFBD@V9,QcI2Y5(\)T1f2YH^QHGZ23K3a
+<.-OC#17(PD-BUeL2e-HF:5P4V2Q7AT2FB2?I5&fLH02D5VW8PV)aKaMP?382TG
AX&>]V<Y8LR]YR+63fLg?NB,QcI,+4&Q;F_fg^g0b#PCd9Z6V+)Wg]OcQ^O)X=^/
d;d3:#2d9N8g[2-^b;5E9bV@)-YO]PM[g;5UNK(41Zd8M)RFV.WI5<JRfDcbP\I_
gS;W5BQf3GVEJ<6Rc:<J,aMCaW0Be)K,VW)4J6d>8N2dA90TLf;AgC9Q:WgZQ+VQ
e_5&Y6&Fg5#M-4[U#&XXZCd/bCOaC_f9(SaTc<TVA,Kc1Y3/85a#5@4?;U)ZVMRU
90D(abI57RbJ25ONUVeE;55ZQ[L5#9\^9Sd82dQd<UL@e,Oa7];^S(UN,3aAS>V-
TLN?f[0gOO,)HGYgX;AS10C[^;)>4R7;K;087e;)_&RYZ<,YTE?PGB5U2;B)OO4;
Y1aGD5:J5:AA.01,A3H1c7;5SXFWdWW3.7G9FWIe,L9O80aXL1=(_9eeKHELGd;]
9AQ1:V;dK<g><fAP8H:/QINVg?66;KK8Z::X^56,Q\/Aa,ZX53Re>Ie;Q7J?H(W]
a_:eOPK>ScGNab^/VLcDN2Xd#U357\-dH18[d[1dfYVOM#>F2d?7MJ1YLfJ\gU96
HO3YHA2ZHRd/e(P6Q/T7NcDdFZ=<Ae?H[2_d7@QTLET<CK;>4.N-Qe_]dSIXKOUB
RKd?9^0;V?CB[XD0Cd0(R486bY-,9Z_X6,<WN;NOb&KJJDNMJ(.F3E0WNBQ2H2@F
a)/daCDc^GVdbX?Z),F#5VZ6Y.V0#-C4D4-f489]DVc3H@&Q-Y5Ug#g9^09c5aJW
MJ_7VU-4e9bCKB:B^@XU+\,0DV=3g;1K.&#-52Ue4fDF_F85V?23(f5b<MFQ.H&Z
Dd+4G@,,3EI<]:RRVV#Df30T)7EO2CBMTVK=L6T\N(NE1\0dL+TfC-?Gd=L-.XV9
L<>J79YL+\PbPO,639N#?YebZY04.UMe\<4>[(g>-T<)gM/J>58_N:9AAS2b6QB4
Vf/(,&<NbEe(@Z&10^]G;((Sb>-:XZ6S#HD>ITJENQ[O&]L?+H1W[W\H^ZE4ef.Y
8QL)c+1[6O6SWgc?^#+L925R7<g:EDNc5ZT4H9DZdcbPPd)\BO=NMR7a^4&?)eff
\d;C&ZL]R\)7NTR_65T9cRWe2PH_^IRbUUVCaJV0A3(W&(HILUc;D[#UdFb7Oe/W
9X7Af/+>2:[EZ@R#D1d^1M5ad34&8FN#-EO6ag9IH7H(9SLBKa_&RP&<E5CPC&fJ
)Ib]+HRX--_XK6QNHM>CXb-UH+@=NYKM\OFQKT(@#7,J1TJ30+V,1#U_7(3IR4&,
>&#f7cIa0aCL-/5(<FYC-3^/\9;JXI9\_+]9+-_aK1./d-QTL\fE<<^##3Na.g@V
9MW2gcQ\/4[IE-V5G+)6\QB/WD6ef#,H()X,2RU5Yc=B:V140I(U<9c41=0,5VL(
W0@@aPg_/\6@SB23FABNE&6+>L^JFa#9LG\<:[M^RBNNJ6+.UO47,N@F6]?]\cfJ
W3GHPN[==R=#gFJX-J2@b?bCI,P,,AfcHJXdM,K?f69]+BA.39P#6U8UdK72f,A:
IT:QE.6.#:?_<EO3&QGG+ZH(5\3L_.F5QdVO7I08aM3HULe)2()2:;afQ&7TNAON
.L@V-a[U+#[=R^e#-@SKVa^;H_I9\GJG/af,b&CC_DU5EIc[))YHQ#eU@H#&UFQY
QZge401__:#GeMcTAIfDM=<E[d5IJJEbV#<3<U>N.<\.O:_DH/&MSe76I6+GgDU/
JA[E)4eCHD-ZZBQ&+:7I6>0?>.]e6]IA.W&eQ(VR8<=D5V7N@Z2SSD,I5XaJ^M<J
]57CF9E?#39^ZGF:e(YG9V(X8e/3;YKBDI+4A1O9]&RKQCQ3T1C]^L6H,ABfQ=ZB
DDHK6XEgffY7)D9VN+D<5.UM8.OS#ED/?d#EL.OcU3[7gJEYB5cLY@R=eWIUPf-/
4eH4&[]D>Z?<5L#LQWREZ@daFJ(a6\_-abgcZ_;V8[M2Z-/H:0^II]LLA:#Q;.F0
e]MY45CFR;3C8M++AL>I<-c]XFF.-_,B.2\fWM?/5IbGcZ,]0B7,TCY4G/M71e39
dHJbVIUafc2V-QGcPABXWX8.f4-]da&9LZ,:#3\A@e6HDI<M+H.KIA=>T/Z;Y^cP
6CQaW.UD=GC5@A5?4\S+bM6B[1U8J:Fc@R<SPHFY)XU<YWO4MO7<^&6TJ:AHOIX?
32DR//M[)OLF0?UJ[-bTWb2RLTW\A<GU,,67DcOE7a(=27HQ#Q8M0(8E__:7>W,P
PF>FR?Gg\?GBJ0.5)K49X(2Nb)G)0^?5)>Y5MNE(&[SDa.,SMCbdP\LG-b@d0T7L
IeH;)3,O16N/fSa8:=>,WVcZM;Q^d_-N33)(Z623bNBdJVbfcP^b8,\Y@R5@M9V?
a.&JT0XI@#1a9XW[aATEYa3SZP;GgdfbE0S7V7:cQ?TAcTe=)#A+-7/dZ;OPaggM
H,TEO+b7K:Y7&^+BWH;9aJfE:\3JQ)3OSC526==6,,&,>>(dYOOJe,g8X3aOTK&4
(57+Bf\]b(3RNVF-6dN9[f5\5;dL75U1,+]Cb55GA?V&=&aQL?CG]9-.B+]UE)0Z
3TC4XUd]/IYPg4#e8OOAPbME\H.c[/_;g&.&JZ9PWWCZ6(a/BK@4;QYX[f&Ma0bH
3M4L5c0V1XF;>UD;cV3d[&4SAG:4a(2)X=dK[d,+/74EbV<XIUB=UgEXcCL0feC7
>a0;0+,=XQ1V[3D.)?d4E/&Y;Q(Ie06VVaXR1N0X8[JIR4N\=KS=.K/IP:/f_T@<
,5?[E:QZL5gBH@[M=Dff/BT74NWOd+P@LB7GZ@B/5;f1O?1UZ&YEOX63E,eTN8^d
G#8@D<gNG,,bJ+eSB?XR_fKc4SK/5>Q;@Z<2AIX_fOOB6afd)f5PI#P/N_8eMe.d
J=:<5W+<+7<+bN31>fJ]f-5\V(??<K/_&P[[Q4-LWe14UIZW>;gcK4Q_T^7S#05P
23R568F31Yg@C@0,S\aSKc<L.Q04U?[.UX9Aa<P#3TO&WO.QOTM,?P=4L=>C_)YH
+cBXZ#GMZ+CJ8HdQ=W9O\2]G;ZP4F<@7ccI&42:@I8343Gd34.ER]>6MDQ)C3PZ\
.gF[Z4]O1P<3R9YB161KEBaEAR5VP1bL0>F=UP=3Z;6/ES65\GQQD8/KYCX)?[8>
KM8bPN=3.H5aP;G9Td]<+L]]NQM)IM/aVO>HEZ/?RS<#]ZV2:(B<ZdOZd)<]LEEa
MJ+Kg\QZ,&W^?(7+,GDcWJ#f[9DXaM/\D^[B[4LTUF=L8;C4+_bLT(b),c+OA-Fe
LB,C/8+.,:e](3eMV@&d,Obce#(^aA43?<R&\9cMP_-Y/0>Zc[2&WJd-e.EL@\b,
_aN_b2:]3aR>@d)a;N\1HZS1Q@-.JUe9=+-(KdDP/73N[L-cP+7GF7S1JLNR+&S]
SDI;^RLP.<9:7]&FSZ>17L<23)R8Z#3Q8S9V^KRT6@ANYWP4]]A(dfHc:0_YCM+(
JbRJQg8BJfS5c-KJK,<K21O7J,DT]EQ>FR.JVE[c4&3:;V)EKNZeEdHZK8X(c:g6
UXE7B+8I7S)bICAb.fUdEYg<c,MS(+3g:faFAJ,@f;C)5Vb_RQE3:#&KD>,4EUE7
B3&[bU#EQ_bf63DY/G;b6HUdE9-:1RHAaD3;DR\0W+MYZec/T^]7O,W&9E5@J7H9
[eECOGK@;<15)f]SHW_V:9>(c9B-[R:W]dW4U-C15<N9@d0,RQK<He0Ve6OBKCDL
B3T7]<N7_6SQ@DQHC^X1ZMM(-57NfHaf4+H:?.cKD-=DE[V^gCA+(f?.T&Q9M.B1
.5BR:d9?MB((^6g,XGUPf0>\D/JPS[M+<7B6-9E2P7fcb_&fLcS.e0#Eg3)4),EC
a,[K97#WG_OPU?MR>P&+=Z#g]RW;5KA>NJRNRc\2D]S[cHAH:+IO((+H+S,+IYN,
ATR(V4Z53;V2g1Y>(:YYBLA-Fegc>(X16ATT/UaF(G-1&86:-#5CbI9PR0#D?eMf
^.)-AeJ8^fK#Z/Ic-/Y)C\Lf^3+X7MD)<SJKWD0WSKVVTOMNJH0JWO&U8-&^b][@
<9:Z;#5P^B@:IT6LcGI=BDc9eL4Rd-]L#IK/P1([&4(HXCIfD8&>6#U1/+ffOW+Q
cY_[<d<6454[bRe&1DO:6G@)_^,H:Z-\LRe)3-/U[?0(NBDcJc3VTUaO,?6WgCB0
+@DPBH?LZ,BPP:D<EL(JOd.fP_SQJ#]]=-3CX@9I\f:I_(PAS<;9:+NY9IE+H;82
a5MV^5+B/Mg)?#e,W\5?[\=V,Q@7TOY=c/R77NG<(J/3XJP<;\/67^:dBdeaVUdF
_f)Z#T?V/83Ec;9YT\AeK27WL;E6BN/XHB+]aM1,>QR7[JI:Tg/BXOWP/\H+H1+c
2NLGe<B1F4EK;+eBD5A6/fE>P/]4e\S37SQNFf&1QbeFVH^>eG+_6Sg13WIa;W=Z
)8Sb8?+AH#57^#.VC4=6)3I6T>^.DfF>U/HAV0SQcVZ).R_CS&3Wa0#48(AK1R@G
.BB<ZcK]6KdTG9]=0b0XF73b-fA0\SaUWG5g[J;#,C:TMC\L_S=&70:=#/];T?<_
/8X:Q.298Z#d9d[/7;DH<--+1A^CS0RcUAZ7:;Q8UI]dLRO.>,ZGE4e](J/+#9Od
#7[))U2b+6FAHKeBM#4e=/1.b,CQN_D,;&KZE[dS]PMdA0G-<FWGJIVM]>4B3<@6
aQW+cQ.5CK?+)LeUe]<Y#&#\3VI)W=BQ;XKOG^Nf(94cPSfQ9MK>_MW\]Q>e,V>.
)gV[8Z/=4OL4CGbK>1>>\Q6Z.4KX15]A^WD=aV-(YO1-63@ON<gDKEK7<\QAKE#[
f])R7-dJSM<L[:YTP5IdE2IV<QM5,I=/>fB]NV8+,8P,b-a\@fU<=DMCD+69e)^^
;ZG6#AH@;:6dMgQ:?,3fG3KO#db/Fc/fFSbXJ)T1e66+e#84DE2H#<e/AYY2K8[[
fe,33?1^HI84ac/aK(1Q/S2:\,.DaN?RagQC9_0VCc6Y)17^OX69H]G=>,5(L4F]
a(#5QH08[gFE3e2N3V<^.[31DQbb^]T2L@SWOVb?Lb7MSH?Q289LI;F5:#2<C#3Z
N^//A9aFX)(<SYQ5OaV[CG#^ST_GBL3;0Eb__YQ;F&feTC=9YTF)F?A\BPM8Z0FY
RK.0,KEY0NAJ++K_\:J:>3HAW0De-,37Q\IT&d&Z9_<&+bOGf#eC@]b>NEbO0JAP
B?E&1L(8[aV/_FDB^_];QUaf53DJ\:O(Q3fScfT]aYSfFU6IUc0>+f.P<)\e75BR
^2U?ZAT=0X<C=1G;9d/6I,_]6]W#]ULee7a7+gcT81=JE\=g]92:/]H2(AQGL1f]
&GBb/&G4>BDSE^>Ge.@Q\I.IU4)-S.aKFeAcTWJN/B<^N]MI>E9@]9,-X,LGJZKe
d+OA__fCE6W@cD[DaJ&F#_F??&RZ-INE@=A]B(]e/L=+e(Mg(7bT\F1C,C7\0a13
)0>GR[KR1eUPZID_-3R4S#/VSbR_d_VB#4Zd_ICLb(P#RPQCV9?YNV&(^LX+_g[<
H\4Z0(]+ME>(9<5\,KITN-A(\N0;;]ABAM\KF^FD3-3H:&9DY<,2fS8@-U=8M@4[
U1)3SaS)QRWUU@?\0^,7=2O<1VXEQTD_R:UV.()ZZOO\eJ+R]F0HD4B9W47O^V;F
TfXAb:>&V?(CNKR8W3LcOd<fMK4<bG=;/M)9QJWJ<ZIN+>/bG??HNV,-6YN66(HI
aI?AfZdT@gH/@0e)\NQg;a:aXZ#2#W9E\EM?#V^BdO_6?[0XPU/RI,=(65QIe_MK
;2C^_cY-@A/=H3#)3HQ?51\baCHF4FaT]U]e\+OD)25+JI>J#][<=QE/8ec?T@>>
X@Dg-SSf>e@1H=M2,FRBfI[-,XHA(+2gf;?:+6DK3\5]/8C(9.1R6VEVZRI>,&8G
E_8C)(XI.DPD5KG<LFEYXb23O8B60R0=AacO)Z#cINQP;./J7IFPdA[Vd2]0+34(
H?N,#9AK?)+,ETD1\c66^U?I_CAR^L2S@.;g)VF/=#d),a@1Je&((\<dC\NU3>ZK
LB.B&[Z^GCL?WY&FOBMZ^D=c)dPZ24FQ>bRK=9RC2O)EKXL^AK9I9BNW:=<YeMSO
dVId\Z=AN=5>HLf,P?7.W5E2#=:R;C_Y0N)Q=B93L,NEd]28)3d^62#1M;IAOcf(
XDU1OfTeHY#:P3A8OW/@J3aZU=J0KRO6G#a.###PEE-^9_c(UF4&H&d,0E=\E3N4
O-#J6<:LQ&#O:7<=P/Q+)CT2<KTe-d;T<c-VN6W2KCQ+\FIH)SGE((H&I(GZ-2,a
S#5#U6B7L?AbKSgS8@[6F[H?ARL96;THQFNQ5+:Oa(DJ#65/9.&OD:HZX#d7B;U6
.1IF85B/9;._>4+W=+-TB@5b>@81W2U\G,+/<e8KA(BL28ROURB+0;FX@W<B&9K(
,>^a4&,2]3]=@/P;N2g6UYCD=B/B1#HMYg_:?6,9)J)eSZ,b6S,U8ZT@CKRNQQQ(
^C#GQ/3bQJ),B9F9f7YFG-@4]S]^30F^.L3+X<WO-e2SQ@I]d@/-RPHL1BQ]aT0M
,e^PAQ_#HYg>7E+9J-N4-X:gBGa)O_E0_fHH\dd(KPYN\X3HO=Y5X-;@f>H#+WA/
UF&]fT/^c)Y@=SU=G1@)T4e4)]a7f:W-:<=#:e[cJ,4.f)bC/8-FTY]aO_f/LTfW
O?44c@W8>4d033&8=Ia&--+[AM225O4\D/+]OABL;?HY)TFHKH1KW032A^CV77UZ
7N]fcDT1^UfOLE80G?:IU_A[4[c,]H1;(C(cKR.\1H7,Y2bA1d[=I3H0XL8]g+a9
P;6J,ecZ=MJ[&>9Y__bfYF+1A]cdZ/Q6)H&V[9^SSXZR8(bN=S1_0gNC:5J?)7/1
gDBU+,a-K-C&R87C5:/gU3FR;A??6C)1,DR^HgT2NS#g;:HX+g=dJC,X&[:cIXM1
Fb<_?]a+\g.gKT]C7A9Q>T;A.CJ[^\YF+^>EP,75.F?2AH3:e:c9<2DILHJ>EXUQ
aHSfGHYY2VC))0I?[?dG16^C9WZ)[OCP^^C,D:>[gL76#GI^<?9N8?NX=d:+83;R
f(M_-<T1+V<TPd4N-V_a5DVa]N8XHNfd[H^#72<SX=,>>2Z-TeUe=<D6+9?V1P.,
;2c&EV@&1g[HMDACY5E]aWCIYP==3IYVBS&;G1c0X+;;&-W]-CPGIF4A19.2-f14
eB?geGR07aBeY<fN3)E:aa(MP2+QJW-HLLa,X&P]YA,d+-U@g<>.NS<QX#2;GZFf
CERZ.E@?659EG7LR&QAbF;6J=E:F6:C]?(P)f2f6b:f@0fGS(-ROcW9I)J()&69,
9G<[+D.OLF)SDWPYQXN3H?eS:=4Y8MA;PJ\8Z,NaCeX79+[=>b@K0=(AD_@S.gYd
g/OFGL[,4=-e5Of,.BHd19bIX?<OG<6A-,O?OXILR?g3B8XEg.8N/<./Ydf6eH+g
2AOT^8Z<;E26=agXOT^Db6cG2W>0L31A\J@+XfI\gB+9bHQ]^[K&42@GBP-fW67b
82Y0,;MF[LQgNG7&);CW/7.EY5P^BT_C(8K)>9\R@/]PFDQ:+CR-M6<VcI<C>#TY
d(fffKJ[8V/4P5T(?Bc9J/a:8.(Q-Kd>-R_K,G9LNC?\JM?Q[/c>ee:YXVHF_&,,
2BbfXd8BX(2>^Z4I@<ILLTaGX_#((3?DHS=c]]5HO?[O3C-DX9K.R1;L(TI:f=V+
JMc,1:E25:Ce+S4?DMGIY+(C,&/PP11Cc8K/(D[)R6.(F.F_Q)1W3-QRR/+YN<6I
\Z6;\=68IFg:(^/G\;^A//U\MfBN6^<?RJ?IcF58gWI_P7NW]WVRbE6EMC)5=\fD
X3U1bD-22<ZKe&HHGG&C9gPTX?GT?feYS,0[WB5#,&X6O@f9PE;O/I[ZcgV6QF9I
J<ZLO,#L^F18b(gLY9]@11K2K7-NA&9L/I=Z;MI[S+58#Jc/H57O#bK?W.X^d@<R
5(L=D9[KC[LR)TdRJa)LH_MOQHe;/Kb2FVH/&G]05#cbPTTf1UW]<>=D4c<A@BS+
5/K9bR_3/@^O(2_:.SIW<-)99L&]=UAJOM<^UW9DF&G(W9AN75-PWPf4fRG8LB&)
cOK>N<[N+&.c]2D26A(>./O/B;5Xd[@a(375=+C39XAK+B7,4?OFNB\>;b___N]]
BJ3aX\K(^?S62>&fMSf8&A_-:aOMU]g_8M>@Z@_NPB[H+.\9F^-#JKV;:.W\6=(#
JP<J0EW,KI+QSR#?Q-MYXDYTE_+R[82O9#9@<JSgL_\KR@^M2d_&GF,76TSA9^5G
A92X,?&@D.AK6L>.<[\ARVQ0D^@1\c;;a&f8Cg4<ef1XgU5ZAHV:Pb3/DI-aL3EA
?a,PYV)&/HU5VECL4Q+Nc@)[5b?g[dNY&D8&dMR9<\2;</5;OW]c5+;V[XB;aL#4
S:\9K;-eO+C#OGD.A?TC07-3fD>VYC4K:)fO^+X;^B>5WY9b2_LT9[4Z&XZ+:/V8
3XKIJ12:W+<(\5<(H61D1A@PM@X[Y,ZLG_=#EQN;7,]gCX8RF19(?>LL>4,aaUSV
MC-Ld#d-1J9;6:9#NQ/NgG\SDG4NO[E=LPS+F]O5,432a;-ZEEEeFOE=AF\+>[5W
@W]G05;,LJK-GIM#:XbFZI\#,#9D>\)3T2(WOc/&&cU>1Y+,@@#PGT\JF#Va;GC(
_)?<,,I&)7FR_@X2BO&0.^\cI49LO92Y4CD7gc#4P/=;K?:^CdU:Z4>DZ^7(W2]6
P/Q+\/Ia01:N/7Z=))R[a^B_,&1,/f\a[0Q>aJ9cXa5[+ec0T1;H:>P5-,O3MW/Q
;ICYX&H<\@2]]1^R;OI@HcWC(b;e43E-5_XCXcP]JTNGd:E;\Zfe_=ANeRG].XTN
=7]FW1ggD2Df-cLa,C1a1?KC5/V0?S[2)cKX:HUG_R>J/\>^)OTVXb6.]OA)Q04E
1<HWc8fZf.dZ[B;5TQ/2\4E&BD8QCU<O<6AeS4RRBZI3-N3BX4eQ9cJU?_HaUVQK
4WLIOE[OTN6K+=AA9I2R8Z<^(+Wa4U^1Z1L06PH7?OU86cX;VKZS(NNg&ZI46d6)
6,5[>B]TMd,6Bfe,@Y#)](G.;CfBW>7(C#P(9RV9D1-REG>>DS(BO?3=/HUDbHE(
5GC1P+Kg9e,gBE=/RM]6U,eGBXWIV/eQS68NU)2<P,Caa+d32a+b9PEe:6A54(]T
.5IY9AR+5;@PgaD6<LH]bbYC=HTdX:DacC<3N_:ZX,cFR:4P8FEP7cSY^5-UUIN9
F(/2T:g9C9<KfP2b5QIAHU7CB&BJ?1ISH[7Q-AD<[L\LI7;ab02:3CL702De3R7>
<K/e5Faa^@WI2,XMDZTTEB.:-VU5[VMLW[(\7\484+,GAH-3YBW[FO+\_O]+Q1EC
Y&(KCOLGdL>geH1OFY>:B^#:[/_7M5-(=RLf79WV+;Y)-TVCUSJCd+QY_-RQ\M2,
e\#CG)g.1(09)U/VJHW>72?H(].[9E\C51Pg4A.J5Q)(^&I>/<N(?-\_Y1]c-=-Q
ZBQM6TFPA4#MFC_e[eTRJE@G+);;I\>g>Q_cIHL(>H1b-_-3FJ?(Ab/#Y8XE\9-,
bRMVBfJ;fQC^V04SKC\IAc_<.2-/?RS@#5#_]KSaWA(LJX[(b/9?ZdYFK:#+4=bZ
EK#L?YHR@PZGA6&VcBOP<[_3IHJ][RGDW?P&><cWU.0_C-U1G+=&9@YS8=dAA4E8
HIbTG8=R_)BQN7V9Te]0I-5T60fJ=7g@:6<NAL3<XC.<R#Q).E5)^+7Gf0F[/3)6
?VHH>b4B<:R-R93ULT[66UKdGL-2WB/e#/1c,+?H3OVHM>\FEY/9e_6A-(TfOS^\
:gH1HR0b@V\G5Bb:FFSd.=#^]\9<R=#0S0#OIcWP^HLYTgHd1b+1RZ8gC=BO-YQ/
_T:9(P7#J9\,K[(?HR<=]KYA5CCdU(;.4\\EQf4M;\,5CX]?C-I,;U@>D,MYBZIK
UG\Z;<XEPM+U9F9e;M<(e1[a]PHf_EL?[aNEaXT057PW.BcQX\QI-J=a2SOYD;VE
+cD[[(;:75=RGA>2e6Y99USeDECG57BU87@]H_8YIZgFKQ;4(PYc\XS-EJ#Q<2\I
6NPXB-.MO4#_2g=.<U_6dT5#aM=\f=VKR?CA\cS<>^OQeA65@HD&cY?ZVV&Sd-H,
XG1d\.MYYNGM<YBMW1]_dbF+)(XXA[2_d[ZOA[J[;E1[f2@48c+&M5B#DZ4YN?PG
R2H)dC56J4[V-gJK8dPf84E((/T@VV<b)P:&1+]fORVZaG;F+[JMB:EbOI;DTg_I
:<+)d7cBT=IBWL&F&KH5IRe;cS73F:Z;4GJF(G>V)F?/8F75JC?RaBGWCd#5bfQ1
6=<]SY)-cA[[3T?3OOL/ba&O(dZ&Q)J-6__@HB<?e9<N6-LDFKD<M(XY[)K<IQI<
d8)Z>_d7,P]_>;B?IRf1/?ETVZPM55Ve)Ne18P07;bHH+b0_O>+MS/X/L1:Ja(dH
HD9/)A0eT[#COdOQDaR+N8be_<Q)H>a5PCaYGH2[U.=Y_ARVFg@9VQ,FK<)#>TaZ
A5<[9S)[9I+XPC52LX&Kd/@:NWN9=GZdP<<4<=\Z?cV:)(]^D+WS>^GT1L_/U<=8
IVU2QCaUFII8-M&ZE=F^A+/2bL@]6EIZ467+R9/5:cMFM]2LIBF.-FC.ZX\O#g@U
^LW[HW>cC4_F<<,ZB/8>R\(DB4=([-,4a>.G6I;+/=-_c,[=]6f+4C35Ic,+8S\V
?aKC0DBI+BI/_9P-^E>)dBU?HO:c5(;)E21QO+L9c&HQ_7/SEDP<F1/];PZEG7<S
WUIB\B;)\40aeCJ(FIWD(4c9_.g]R@?e#(,(C\RPZWb@F/D5K-F,;&;+[0^JW)8M
INTdgJRGg8G:9f?RT2B4AT]7@f4)AX7),a;7D&5.&+e6/4b&I;W<?g1TgbLGe@=K
FQAVOW>)+F4@&b-FCfRNR382FO7\WQgO7KGa@^2/99HE-P#);d3CaaKbTG4^<aNR
JP;]eBC\YRPZac&KaU.\Fa7Id)73>ZN,WLKQSJNH1]Y3I=dVDc+_-+,QEgb]KN?]
PV1R;)&b<-deIG-JK:PB7-NH7YK&b?cW\(46T25+G[@&X9eO5Y6VCBU2-b14,c?c
#@]QY([]\_IWAA,D<_+WT#[P)WP6FRIU&<f==DIHX\X3(a.Y&=IgV()Y-;5_LUOC
O?;AbR)R_)3GN^S0<Za\U=_R^>Z9G5?GaPTF3Z;M?/E7W3GJ3_CAIAU2H.AgI\,I
D0XH@DS11cd_Y9]0Rc4IcC@^UXLe_=Z&J;KbD2T]+@7K[[cMg98Z<>>eRH=W0fST
,eVSBI9:X@)W?Q>FfTY5766M(FB&7X8EWC[cE@0[YWVY.c>;+GIKgaZ80VNSRW2]
D_BXOW0A,UaYI0I+WF_S_(>YF@:531_YV.K9@I?#>)3=0Uc-Xc_2@T(OI/PBTIDB
&4eT(213^JK6-ATK6.U[.g#>Uf[@YNbKXCZ1&d]-fIYNVMLUT4M9L(e[IA]U8Q/c
/S.#BU]DA+_,G1N(1BY:81F0SJWeFSC>G-^0+\]G0<O]1ZAbYg)Dc;6+]1[M#2f[
YTZ#b?,#+4[Qd4X(=R<T#[,,5#57_VORLgPDZLf7MSKC.AdDG]+,Z##eaT:+3aGB
EO1A3U-3ZB\Z4eZL(9MX?[C26J_#(+6?9^BRf:18.[7/5A@/#7eXCEJ0beE5]+.+
/>Efc,c3#b-1D:MA1LM=H1L5=/]FI0?F#G(;S8L-R/[fT8]+dHTF)E>?^=H44BOT
]@>aaEX?#[5.5+._]aWJJ6d./d?]5CYW3,[HLbG(BX-@,X7HVPE@8MUZ)MF=8O:C
Qa?/L+4D>E1aX<#M68Hd9O+aX+QM2+H#S()1EAA?GM63E5PO=L#5gI?B9SUgdW,<
-DYOM1bG2Oe,:>Y+95\<\dV+OF6dS1(YJ=JH?OX]47VAc->2\Vc7H9+#?Q_GaR=H
H+e4R\@=_H/4Ue4gG.K=&RNUE\,c[;?J-7c6C\I=Gd8P^T3DaH[Z2AXAWER4E[:/
:\E>YJU)6(]ZEH;>8Pc:e,L7)P^QR61QOYSd6/Ic)Y75KG@J)aHH^<D-(@b4KJ<@
/^WT#7QdI+T<)XCCZDU5F]^FY6:XdJ^O.MLJJAYeYBBM@(9^F4U7(0#WW3]e+;A:
K/O=P#(aXU.S8>\Q;RE\cOEQ+1>(B\&OKLHGJB?A:-D8Zd.ARLBQ/VV22G78=/Pa
S2U?[ZFC(TNUV.-Ra+J1HAMCO_K-[DTM+J;B/&.gNGY];VN,@/X^?d.TPb-T3RI;
[-MTKJM2g@>]-H&65#T1PY,>H34dH3?8+BAQA19E+&#VM#C;//1cG<N/_R>5,+Q-
P;)+<UQD+;CV@8,T=GWFN[BAKDcM+a+1c,>J/N:6I,3ae^MgdE[W/0,=Be?gc.AJ
A)&/FMc3dB<gS:9dae@8B=:NTLJU_#QU@2GO>G^RJ>LZbS5.718PKgeg,bK\I-Z9
W:^7=RNN^)9OGecf?E#]<G41@Z@;c9FISXN&XPOPO<(YEV8(CL=3c--8EV>J,6&_
2]J<6LQZI::9f0PdAECFL[gEf_deLR^I#X1&HQ-@,5Q7>EFW2,9PE,O@+I(e@4;6
=d(2.Qb06::/2YTa.fAMBB@0;-,K?PL9,e0GNSdc(AE>([X+#X;[DeN9Cb[980e1
c,fe>]88I:^I69<:GQ/93LK?d+JL:XF2-KN(BWYS0d7+.FF;@[R9J_cY[&Z2[?^U
dV0M-H]T8aL\_+=28N5S&/6S5]N9/X#aOb-878VCKD]]U1>c6?[@PH&D41#I>9[\
G4&YG)JFgB.7:6ZU;9RQ>Kd55Y_;LVM7gMb(QJeJZ(.\-Cd4G?7bJ37K.eTM+;JC
IPT4V7MfC<R?5gbU/Y^B.<dPf)EKLQ#\^UUd?WM0N=\VDBG6@]_2eS5W^NM2GE:Q
[@GRIbW.71E6HWN.B&RE;?0W?Y<X---\:#&eES87IEK^EcV0GG7H4C>?d1_Z[4_\
c:G2#6<:047,7SXBW_eOf91[,#)XZ04AR(9:Z>,<<2.\gXB+If(<OFJ<-g>@73c8
RH0=-G#0MJ+6[=5MRRE_.T&+1D.RRc4=b?d=_G>g/R=M9_WMeMP4:.dBM):#QYU+
@UN@/.B\dF)LU&WDYI.\CZE,=\GP9,a3^^:@X5=D/Z:<L?8ICICXc+)5ZCe@9>Z4
?CI:KIc]?I#NX1=+/8_62a];GaG+,agQK?^8GI9X.;a#aBZ;Gb(8M9KRX.4bI?GG
(P(PSNCb<,@S<S?N17N.WXIT9K[?HG#Bg4WJVCZ-?WK]PZXK4R=QgZ.6#J\GQ>_(
Y9g1AMZ@,J/Bf6M>HMKR)WTST[I8#WEVab03VF\IFO?/9OOQU;F<FS-.SD4P>L11
&BI;MB=UG=aQW4e#GP&M58?+5;SJb0H67>\b,5B+<RR?-TV3W?3egIKTFT2TIVV?
-\M?D)&C=;U?#ZPbSY5:b0Q/&@e_B=T9)/:C2S#SP7EaP_;Q4)Sb(=7)6AZ9/#P6
;W=V.EXSf+I^OCc8)\M9^>UX@Y>I89@X]G2<4P2:-?QB;Z69RN@WQ<&K=VP\MU6N
P4^V#B]B\IW]R0F);a1S)19a-TO\O1.]#0Ka]\K#a\NNA<dGU>:WPB\K?U=J36\6
,K,U?;0.EM6F+7)g1JH,_SN5H<FM+A\3]0eZ.2WBNTQ-4bD_2&L=^d[JcE<6HL].
[.^QfVL^;4)PDS:)3]7P<6)AE:#fG?U:N3a(LUa??>e]7MgZZg80bf\Zf&.>76@3
@f/:fFZ:(IGAA7?=IHR4KL<FUOFQFXZ4.SfJ:,91LW@D4De4AV1,HgX8^dMUHEPd
N3--<J\NTH-[K#feP4X@ag.cYO+MdQV8b#.A;7I06I@A]YEN;+SG67)@gC<,R6O>
XQ)OWS[LGebW.f)/;gS&XD4-WNSJfT8G#,PK@Mec=XbK(dLSFP=B/CPEI5MS@_#.
>;<)^L=RVA+:S0E/#.5PH5=cQS,B391M6O2#0+S4/>g,/E)c/4aE3^)VNd.T;:E-
3f;bB76T+C(ZMObTFR7T)H]>4LXW;f+F:e0DSb]K0R#Ta<L/^(a,FKR;?eX.f9Y8
^-&4OWM@]Na34f,4_[R/BcY4?4]4(_C=9c;Y90)WSWPJAc1U\/D#aEIHTZ/T@8Uf
9>E<YG+7A3<4R;Q+[O2YET]D:c+X+YeF#a+Y]cgKA(/e1]IDA,YBPb[;=#FED)\V
I;HY.NTMFXQGD>&:b[C_.a\@XK=aHZRLS7BVE6HC[VZ/,Y3]A5PKPHd4gCV++W_M
#8,30SXH<8Ke6OPO/Mg6(H[P\:]T9=[0/VPY3^[ef.;UU>O(UU(03O3N5fOb1&B5
+]XSf)T+g5R.1A2c2RbUM0/8R#S_U-RN]LSVX^WF#\J@^X9]MIaEDQ[:N4))e&ZJ
aS<8e13@E/7;eY<=\IIgF=cODfD4Z@7Z>]M<MY^c-C06/e-5AR9.g2-XC^^\P;;[
^YYQdgW<U@(30Y7(USZfd#N94>Tb<2Y0MQ0,dV6aJ:SA<Z4+Q;7=O9fd&R;IT;@#
^\J+KOdQYNS3\M#bc:eEdLUJ[[#gQ[9;C8ER;@0)HR^e8f#1@>NX^ERWHT6ZcRH1
WHM4^HD[Kd<GQWJ/OKQVN;(e)HM92P:P:_T_E@RGX_/2_<g9DW^HO^Z_WFO7V9WL
,F=(EbHP\NXJDUVZL7>GX#89MSKWdM1WJH/#A?SQAf<O7<OVeVE,5LS.NTB@9@+K
R21O1G.eCR_]W#QRN&KGPO+7W<?g)XE1c,?&AQ:1F-&7(,++,^Fc;GK(9d2[Gca#
KQ@;cWS<R4M7/J56cbTg0.7PP_/UH&R3N#76CM&T.Ea+:(GY&0\\1A&<U8M+MC&)
PMJfAV)E\6XNQZ<Y5UTM8[3HV?+]&[R1>/Z1K-;OOdY[@2UUQ\VYNBf.,H:=U8J[
:D^<gC)L-V_afXa/1@Z68@#UXYW6_UU1,)?\BEEY_,^C,#+JCP0SN(bZAI;<U/UU
CTMDa(,/,852?I/87_Sf38KM)^f<P\gJWDNS5g0294f_e0b_PW&R^(]&]O@1[X9.
gWTc.e\4)PD_D?GC,YbK9Y_B;Z8D)cJ/4Nf#(Z\9bGW[DcA:b)77IGgP.8S4,@@O
2O>acc?4a5fD@>L+g_XR9PI<P&(a_8d(2.O88MTMT8YYgA+BCV80D6P@DTVeOWLI
YE]b]Ed0+19172+VJF]A_&VV]d?H.EQ^^C&C]TD89.5bbE(BY>R9:E/a;dc-4X;H
dB>+>7Q_I(Z\fOD-/<M79=,Y7UO-IRKRAYec<F)f&F06+3F>dA<(dQ\KeA+1e0a6
)Y>UQ=RBN^?;QTf#.Z0aKS&K(\DEc3J7QV8;^DLN>9_]X5aDS,(;E--RD]/>]7S#
<YVI:107WaEO]]J))L+-=78S]cDMMA66RGJ,YJP4RK#JY?;])W37;7H@cd=,__1\
.b\3[-GC0D^85fWNfP(S#?8H3.bM5OWN>g<g^..+GHQ_]S8A3@6b_2@AO(Yd[#YG
07(4<((>=&&;L8=3X_1adL^,;[f&WR(5LNFARALeg0_M(M+O]A#;Y&8MfQD42C5H
Rc5cWXQ=1MW]BQ^[=YGgM<G4I>WI(LCBFAM4GBH=>-PVFBP;B/4fQdR86d.b,XQg
&Y+CB,bdgJ:RUAa(T<XG4W\.(Ib-eW>)/C^QMSZ@@#Gc[bd/48Ud=:cM)\LLJA[C
>?J3^Xe.#3MF585L,&QFE\^=)7BCB>A[DB@]V/X_f3SYRHRJ9ZF#I99UAT--R5I(
I+>RNL6Z3JZJ;VLPZ6.;8\3UGDZ(#]c+[ELUg/TfH#46A5[?OfAeP:-WMc@M+N6G
T<4_\H5T]8(aZ-N9+<-KSW<H&ITFD/L98ZfH45VD5,(ZaU\[1cS+7gcZ<XN9H)-^
fZ;5/OaKCE0d+8S.7E\F]U(3c<GQC--+Y;e]PBVV;c?DL:X8^L039T=?7e6WJ:F&
.C]9@2W\\\5cIPSW,@5g<8[Jc1L39g+9/L)C9_DX>(0/fCV,6XL@;e(,3FX?c7^-
PcZ#3?.3884DKJaae]9T+^NL:D6G^)N_e@0@#ICEf=4C;/#;E:BHCN(0YDX^,,L\
A[HPWfRVfX[P63U@,dU.6ScSSg7@:W=A-A9V&JfG[52Z,>^)ae@P(:bF/SSHSdE4
V&N;9f#GeJD<&YB-5LBT3Dd62&WW,A<g<,DgCDD4V7=#A]HaSIN>RAc1G=.,XSH5
^V8C\XD-=4,ECNUJgJ/bCQMRSDd/U@>1;?S4WZZ\3Y&NU))LQY&@fBU;EcP/DgLY
Q76#Z^Y,#@N.cf1dAc8LC:GTb4SUL(3L4OA89d@@27]4Oe[XYL+_\J+1?<H0M0?&
-WR[a<,?>Qa/_4(<\&I>UI37_<-N[\5<dNM63a-@]Zc]?7&D8g@81?c1<5_D#)/b
R[X?>D7fQ5LJc^6e4^QO(USXU<bKg,H/MC#Y/(4\O9YZ#\I@1X(F1;+7T5BZT#L&
6eX+HUZ\F=g4KVPZ)c3e1N)F:F.Za_M@J.:T0@7-eRa5FJ^)fOW521LCe\eYNaH_
0((_\>;AMOS63/Qa&K1/A3@26aA=eZ;V#f+=g+VYd<&=eY)=6:PC(G6eBcI<YH2,
Ib+SGQdf?W-bVLI57dN2fZ1M<;VQD]OODH0[^XRM,UC;1c[Z9W@QE)>)=6++12cQ
/-FA\a)A[Lc)UM15?.MdAO+E)M#9a&51D<[B]-KG6JDW3DV(3@;HB8[#Y-MV+G#&
\+<R.C2fFe^,J]4VO3MW-8Y3OORU[SgQa[)I,4Ba[^(O25fa0J3KdNAKZ_:9B,-4
1EI0S[GNA5Bcff\&\X<Xa9B7NQOJ:CT[)WW?2K7aW@cR+#,4[MOFdL0Ke9\4C>VH
N@S/Xcb-Qbg(0,a+8VO2RC,aY)E,9#:eZ7F.CWB:_^X7,deffKd)U4]GQUD\^cSY
IIg:R&=XGe:G:]ZVe5,OH04ZZdAW[^eTGIHW<-G)_E]3_B\?08Jc6dQ^Nf6I5>R[
N]1#U2HVNX6?<^T1E.a^N^)Ybc8W<b39I?V5bXdWK4AK\KXS3K7GVAdNX6VWR)d0
ZTU;119Oc_[e?)@J?(?GgWY)EHf])X#:ZJJH0_;M_[Og1-Y3S\6#,[XYX@Cg8LQM
gb2X+:3:BIc5E9dTIWZVN.<d(DTF\58SU&NC)DBKJ3W&4U_,SVCKd>IB/4O)&Nb)
4?A[ASc^VN:LB&.cE-.8F9CG(J3BFdIK.WN?bd-A\K#FF#FR\)7e,03(:6K.?(+T
F^:AKC-a\J5NH6FTHLMddU4bN6LegQ1aOJ3>ae;REWJdG8dd)M.g>Zc>.(R(XQJ2
@FJCaG@@_QOdFX/OSJ??E1CS.O&J+33fYHf(0B3^1#KV&[)a2ed]RFU#cgS:XMK-
(NF3baZe[5Q9e9F2?5OG^Te=G+Qc6^Bg:RV9#_bQeR@BG\\EW&,;XF8]&J^)RU36
+4VN<\7Q]Z?RX^Jc_AV)U@;b)eR&/Y>V6TZSb+VM0L[TQ<;L(/7=-0.ZW8_8_JTI
RK8VYdQ];#8U>B;[a]:gC)3Y&,\YFOLPJ9=C-^)K2MT+U@0dD1(_b2SLbEU<GB@:
SX1-3].eXG>QM._a16]\6Rb&^18MD>(R2PP5f5V97I3a#?/+Z0@>71MWQ[CLaC;d
DJV61=._0;O=I;0/Q#1>IUVAQLe6AW>OIF-BC@3#\U0Y-.3LaK,J,fQ4ZcN>:ac[
=FI/JBXR4NdO[>-UP/\^-IX9E[WRb&O-YOH9NF)+0[PL+FCP)F\.\9L\da=].R]3
N>Cc>M-YQ_8#:?RS?J24-8G/d9d[P(5M+:^IWAHXF@QM&-H<A,gN=<3dRLfTQLWL
eQ?B^WE.G>=8CcJ3OA4U:TG,cMU_EH[(?<QI@?L>746XV/@+HUEW\HEG/?]TI3Pc
+f2@DARRH2NbA4G@+CFY(^e-F>/QZD>AcW=3/R0Tf^\]6dE<QJaA2,H_P0;LF_K?
#JT&]VK6;_fEDTT@I[8()[;?P+IHN=J5[@W(9fK2[O+.SI1P\7T923U>?HH:G#f7
Ibf9Z]E&[f#679MO^>c^/:1d\eUN>_2X;C@,T.8SP49&YP_AOQN=f0AB&2[1bc=R
^I<IS+70>:?b&b\FA2E==[]U6G/TMeM04BPD8BMOTN(&,30a=_C\+2D75</,9bE@
LgI76XD)P2P(EeCY0=Le0=Qg8U,B(I[,-2=_2<AT8[:R\TF8TDUg(Ca4()6GRWK1
f6e6QX9TR>GA\;@Z@a4#IaE_S#]7NcR^c?T(3^E>DLL=dPa0A1PaDG0A?YEWP:D\
IYI+&RUC&3&Jc[b2W6QGP=RK(?RLV[A2_3;>51/JEF/f4F1C1WS=]7Oa1:&fK^A)
8D@:W0V;;V:7C[]5@A-RZ0(:?Lf)>21gC,).PKdKQB-gFD^^[]3UVSRWFRa21g@1
58/]4Z,6KYNd24]S#]X@UUO_<;S8QZ\56ZQIWJ.#:G]^OJCG(#WcKG.;g0H68JdD
EK.PfF3^MdJHagS^fRA[PCU/7_,C#&)Te>e]P&@Bb46A>e(2b/DVYDS/HMD_]A;]
PcGcaBK#eNH.^6-:_;?[>LJ&J^]Ua-d4eb6PSG?^A_+W+82WE9ZgRf6B9(5Aa5,/
ecH;gN6Z+?K<-AeAe=5He]SG<MQM-Ye((G=);RAKT_SRea@)UP&3WOfU<WCHHBS<
R1eM4RN[SP=,SKS(#<<\O(ZPC5:^IXa@X9?BA1IC)A3U7U)_d6&=<E]7IM_FQ,D9
C9fF4@C;@BC0@R1YP+Q>64A0+G>f/SS^(RMKE]B[f>87LW2.CG:;E:(^1A&:Z=d&
H:#\#(D0/A5]b>a1bFd,=P2K2IMH4Cc0fI5=>>)Z?PO2^H&/aFWQ&E_:XSTIGX63
UK]8P6b;07:9a;Yd)U;4<\#f?c<KaRc8X<gf<Lf:X)6Kd>(OP/g_CR)K_?E-<PX<
Z0Fd5N2^)_gdD9^UY7e,[_7PG18gb1#A2P[8PI;PQLPMEZ+4WED5-MM3W,7(XE#H
N0?_5]WEU:+OMfJF<OF5TI[]c46DLZ7/I1CXPRCV0B9.6KI_T1?8#Ef5U(Db.8=J
[fIJ0]-^=<2E8);(&MQ,0W+H\b#BMB7dKKXV4MgR-@C&\f_VOb@QU)eS(O,+UN+e
KY>:8M+39eZ#&NOYV,bC<58>&ONUZXL[8JaD&CKS>e=:+5&ePVP&GP8/Y[(V/GeA
>>/(7fCY/7;deZJV&ZF&.AJ93L8YU_II4Q,gLMd[AbfgRF6BQec]1/-R1#82Df&U
.-RS/GC1W[WH,4THLE^YU7aUVZD>3=bA/RA9<CT1WI7(I6&&RO))\Z<b+RS)(gf5
g;9Y?@_H(Q_A5P[L8C1Y5^N-[#b[e3FXZMI.<B?8fDP6XTI,#>RFJ3A4E]0])J@+
)d-W6@@J)\.U=:d(CWNXT;FVC90AYHZ<CgO4]I\fCZ37&U.OTd3+-9M4JQ\DSfD/
QU&PNQOJ9OL@KCDK1\F9b=QO5QXWa+6L+C7M[;<ga/a?^]?[4YH??R\:+PSf9TJD
\4IP\&)6=G4X_@AJEC1K+&LET998-ROL[Q8[/5+?M<]S\+F8:&^H,61,1U2DgK4,
#1(PT6QGge@4I[)T>7?,_PI)_]:_IODPTbOgI/CFT4cZ5a@,1],Z.,.4?QB#5<,@
FH<?A#.g-6_7a/fHMR7[6T0_YZ&):=N0[g>VNUUGf+R_RW8#@Y2GP]Pg6W#AU;gd
TL4;5LS-KNEA\g\32QL;H7:JQ9MRg(Z1=&-J^I#Vb1J,]\2JA]>^e]6PYDI)1()Z
Bf)F-JH]=EUbT?9/MeT1OQ]6Q,#BaO3bAb/6]<M)MH<eB()0G4@XZS54(@a8bL#K
\bJVCR69IW9R;PB567IXfC+5d8^X\LDPQ6S:FgOMbY=<FL)^M6EN6/4+>5FB9_F#
K(^7I21(TWZe:^;_S;2_,EU=-TbKXMQ,+BPL)9HTR:HMCF5,N,#J#V8.dP/C1>]-
Y-.J+SN/+UbB:RF]QCgH-=J0N\5?)^)1[IYUESaa3C3J_gM1;MeJDXIGS:0GK:gD
3O#7^FU=Y8^O+&f/b#_31<EcEP>3Ja_/[_LCD._WBG;-XFBP(AQD\M/6RB6A4U#c
)JG^:^H_f&+(5Y#XLE)<O4+cR/0L-COQ4?L3?7C\Ha=O?a389[BO5H,V\7>(?NS+
+5[3\_9O/L4&a,O;6K&RA.B9449\&)RdY8@_)J(_]PCP1WS@eZdMC51>[#13b7#K
>G[BWVZ,,AX:D7YL2P5@)3H8:R?X0>AU<9&_73ZPe[g-_EVe=?GVNNF(HXH<JeU0
]K_dV:G;,D^JG44_>9?7XeIUJ2cd7^PBUEHMcL>,G]P5^2D#a4VOR[)&D43N384:
-=UQ_cJ3Y#6+ZAABbLg)8ZZ>RZN6#(Y:/?e>\&[I5#7E@:>&^^/M?a?&b_Kc7FR(
^Ta.17Ac+3FE9OS:R1927Q-2[2##F4DRT-fG-V,(-ES8Wf063RLT@,83+5OS-7&1
<-Q-.C1-BZC6=>cgG>e5WRSg><^-P>_4YSH^V9>(SbYB3P(dNZ^PC9#0FNMG:a6N
Db57PLAM:FYHXb<+Yg>;[88YMdb=7/cN[(d2c4g?KIZ6F[:52BZ^5KGE.)6?:X\W
2f=YaM]Lc?&RI59PA84&06Id@/Da_)XAT(^_@NT15SQ8&FI\6)88b794aWd[ca(5
fF/geA\@\A\/HUVgIbg&GA_XAB,R,I/>Q:.@H+)JJ:M>9[J\G>=@9SZXDgC(7+CZ
A(aI193eSE<WW>7]b&>H<4L[<2-Q<K-\&J;#(7C=bEIYOa?c6-DV,:@@7e](3@?Y
A_.>e]LT6G,:JGUQ4(P\.4)/Y(SR1E_D#SPW0TX90D3K[7Y>Z1=LYV_5F^(]YPBL
O_7WG+(O#?1a_.SFa(BQF_5TfC>>919LB0^?@04HC#D@[SE6.HA?#5g41RAN;e;-
NG..SdL:;<9<;Q.KC.8TeU<+fcCe@W,=^O+-B=ID43OPSOAgI9;WW]K5WW\NPMH4
^0/UcBdM48HW_6Gb[48\Jd&^WJ@Wb5#Y,USR[a>Q4E+_B[#>\ZH1;8SVA/IQ6<E]
)4N]#fRS1,MH+Z+?-Kg2+G;^Oa8b.;2G9&1b+cc@Mb;<FVGeY.6[cW_&&Ra]+06g
bZ4>=B_SF:DF^\K;-4c:2]@J(0/M_b0#;EIg:ba];Gg372f(JI[,b.#-A\6eZc[K
e.\0]3Xf<AAGN_MFR-E]TZA#B?1G.?_9[=C8K,?/SNG:0#IF53cN<_Id&&I)8f..
^E7@+KW>0NA\_.41VRDH5e=4]5<@a(<DLUTf1@5TX&>&]OYFY,.O>RXD4=KV2B^)
V\EE=]/Q+PVQ[FY222dQH)AA:fE/2<WG]SA6fW#JN[#V><Y.;@P;gb>>J1QD30b&
U<-:27Ta9a?f&Z2@_YeCgC^J6#UHMdLLG&eePW+W^XB@<X3M(9EgWBY228OX9f0P
\?/R<Dcg6D7UK).P[^MK@dWD3ef0R>2CM),RA.f\cfH68;>N,B8H.(R(Rg@[eBR)
5C:-Y^A.FDGXPZ-OO[c;7gE/#3H[:Ke/(OAb2+gTb5T?bI;d/K6/CR@7P33R[YVC
3>0C0)G1bGL2B)c#&A7;JgDdP_Z17Y3@eBXLH07#Z1aPd[B[NX,8Ke?C96Y.=1Ne
,4adD5_86NP20AG9A33U([X2WHcSP(;/L:fC)H8:=X^PUZJM?#4<V>U4?#KV>AVR
T]Q<B<E_@?;^Z@AIeQ\3ZD<A,7.Nb>^fLL[^daB3]0a#M3[/\H3B7(CA.^UT-6b7
TEDgRA=/NOJS9QN/8AddA.-.L\eb0feFN6?N,)[Vc5@@AB/<QdW^<K3?JGD+YJO;
5&GKP>I1)d^cTaM[L,I;JGVDUQ7II_D,^/1BcQW[&\QCgfA4.[^8^[E3T6A,P[LP
_07c_Sc:.[RMV5.#eV<^eMDde.G)C17)S7McPW6JgeK;X)(1?X&J/@O7[=F6BD\9
:DC/6+@I-GSN\XG/,<ICC;U>=>g+\4EKYVW>a(dTdY1;6dRU^J68MSNB+S4QZCG[
\8Ha@.K]&WgedMLF;,W9a/L-,N9PO^7^cdXW_XfP=NW8I1Mf>eQ\R0EJ)^N@UI,@
_?XUdQUNLJEG6Q0O-UHCYIe000-QaSU1C[,/T^6gY;(?A\aNBG1ODJA;X=Y\A4A+
^88f(I[L8<=ZX#_f:,I0PWVK\gcf&1I6e:V0]ZK>>[f84_?>?-FTE+N5#WZL.fEM
O88;O,FbP4a6D:^ae6AUGOVFC/fLXW]FBDE.(V6HTBaVP^U8O1UF-VOM7)D/L9Bd
LU/]<aCNe.K@cL_=YVMUTO9)4ULEYWK#c0;]I8WQJdg4e^+<KLM(/0B#QBYQ5_4-
FXJ@_0=Z0##-=)24_>;3:XVLZS.D<V)-+S?aU\gBT6[:d-XF^AWXD<L3-N1^V7FE
f?:C\C4YDMKE#VaJWD4[c@4fcD&OPD8F6Gcg1.Q.cUX3F3#X5fOaRSJ_U)S,4bNE
+0WI_;_aN\(7<@EfSKTF<b#.IfOeWR2D626IYZc/7D__4X)>S4RH(g<BV9a&W1C@
ECEQF(>fL1b==[>@4L]2.6TCd[U9,[((W4cL_MfQ&G4<N(8?)b:^SgdN:=g[EcRV
;b4WCeBD__D>;4cM>DE(<7O-FV?9C?.L2)e&;&IK4YN_G\NG3BLgbeEO3R?=gBN]
LOM))55@WINe_\AFPdBCL0&]f_S;;;Ba.9_7MOV>DPcTL<O[4.FI8USH2=?/R<JP
(cF2))gAK92ef6>B;(FKCFD861N]Dd=0VF#K3D714XKaH2W=YF<?.9b_M0E2V_HZ
UMIe4N&L_;=^e<RX#>R@OM36?8CO6J)S1P.@5P/+9&:E,[/1VR&.SN(WbT6CQgQa
^8-3>]V]gWb\OL]B\IOefAGU10B@/A8B0J+e>13g@dGa),@#E_/cf5HJBGK^c1]5
@f5CP/:22aGBPKI5Hd?H=N7.-.T6XQM_2-FH\4Hd@1OF,D^S#[7BBK\>A)8E>bJ<
YNE2U8,PGK.F02C0/dAEc^2(_HOGTX<T81BeK<Gg][?_MXDWOV&&/@d]35G^da8c
c989@C1BeX5YbG3S9dF[11?(\Kb;+7P2/G>)BACCMd1)]Z4Q3]NDb6:G>+(Z#gVN
TDU4NGZR+H3I>_+/3g8G9>5e=Z[a0(<S1F=8Zg1EMcJO@g3=(?F??KeM;V?(SY:a
JFIUDU01\#QGf]fF/c5Qc77+=3,N_d0?(\;<B1)]]<:U#&d.)Y#bPA_@DY_BU?6d
OFZC_\DcQGC34J=Tf3C)SX>Q\NJYJ\@EN&G>Oe1e.Rb7aYPB(1LFX:@^.OK.0N:8
9_(5HI\K7&R?H3OF(<&QNf#45OTHM(OP#<WGfP>&)6dW[b0UUR7TgZGZWU6e<:ZL
I58W9LdE,B6ZMbXI86:TdS>)\XI9WRGc-<1Z&4_EK^E0&P@RN12<8?H(3aKYL^_c
^O6LK#XcRLbQ/16M_Z8bJIV<g@;[Je=^<[OdU2B)CK9<^+:HC(,?BHS.Ef.Ig/D=
?9d-gB9UV@O]6?SF#fGgbC9@:RbZSW32-(dH1T?KGW0BIB,-SI?L[-G/d3E<e8AT
)GKZ?6d/PE5;=Ef7B+81@bT(4/?5LI.8(JDVFf?8-8-8V>=CMHFO)KL=:NAR=][a
PXDN+gJS;0>;T:/L&bKc6MR,WCBT<L8NYP-.F#JN1b6XUE=&ba>fdR;X.ccIM8;]
MX<GDM.U[+U4#W:<W&H6Q[+I&XIU>1/6@=1^D2ZGIXg\H=7]/8d-+G:\e^0E>J3;
]E1:[M6A1G(,ZINQZ,6VG/^Q,XXBRXKY=#d]);c.GC^&.9bTFfZ<GN>O&egYgbM;
2TSD6J?DDB2>8VT:7]9EJ:K3-8:8e;5<QOB=0LTHEeCLKU)KF-&dPaeT)VH5:J?f
C_(@2bJ01Z2MgL;UEQCc:]a(C_O0)(1DY)a+[EYH77aEC&>Ma]7Ja=\\NWfRPV3M
-4@CPJ[1Y-8S+HQ0bfVZ6NdD.D:2dM_Fe7L#\b(aPS,RT=M>ORK)>DPC\I5Z(QTK
B,H0RdgA@6TA9AN6B5WRVCOaBAd^b(cB(5/Lc_I[NCYS]@]f<]Rc\5QJ;:+#^1Hc
7NHG]H7=)PACVRX]T:6@ag4042aJg9:SWNB(-S^K^A?R_MPY<dS,X,F?4W]KAD]I
0]d1LU0<,5WKNCa)&e,OTY&S&&ENLR^AOM;&0]FdHe@XGa;1d5+4\>W^_AR:>&Kb
AZ]1/_WFGW_adY[b6QJ]XggKY_8_FTe]M<;0]dSJWGK[d+?GSD?ZbP;;B=1./Pb]
aNOC2bD3-M=N9fHc4e\BZMC9;57MH(Va@cNdc/E+&H\F8XUE&I+=P:aQa<bO;:<d
Y(I5eg.5E<g5;H:^8==Z2.&2\ELMcbD;_beTeHKYZ5>PW;:(fQ>.^<.Fg<N45WFD
>cU4cHW<3Q->4La9Cc:.bM9L0BA_004cgSgMW[@V>O08Kd,1&,_EJI@0bX68CS]U
8=F8&F<0W2:>K2C6MYIH9\Te.>>#R03LS[>[PCP&a-[:D#-2VMAEVd+&XEW:).[,
J&](CSFNe^aN4D33.@gV57g?S,PgX&gcVK&D6YM(45Ma]=>HUF@e)7C5VUZ)Pd]D
B?UY==[XC#O\Ae((7EQ=S./\:&c1FW-]JJ8#EN?5Y5\,X&?ecT]TK315AKMG<LTV
LgHY3&_?5HBegI<94\&c-YY2EgUJMcUL94MG>\5f3>S]IAP9DKG5<DMK_2DL?^&d
,RQg2gE&PS,4=?VfQCDM?\:D/CELHd2EdP(6Q_Aeg+>/Of8R4Z_d\/GPX3R,(fHD
\WQ4^O:?cUdgB4JAN56A3&T9]X]66CJK8YDBN61/)Sa]?G8eAgbb+<SVF40f9^3T
Ia.[JPN46?\RR14(W4Q5gV@@7N_4R8-Y3<0:ORVO\JU;0=107/=J_Q&HCcMZ[W/:
cFD58ac0QS?aD@HW,U]B&A9g>_0TSF_bE[WYO3FVcP3:N5fQTQ#LHbH..TfMBb](
E3VU-D]+CKQGVK_QfZ/D[1T]KS>4;X3U)?+7).eO<-B5RART(#5UbYDKD7132_0K
+S<&;BFOD03]K&Ig)N-RS+R=.:M\O?X=,6-P_PXNAWbW.9]9CVR(MO)KL^CFNE7=
&+E6CaMX_B+@]f;3_MT+bT2Uc3\7IB3PcUFVMS@Vg[M:e+Uda=^0R_FCQK)P=Y8)
F[.R2MB)BVP@K>RI,Pg15A&N,[453aaPXg<:Ec^J;?Nb=VP=:@39/eW4[08E2Y56
C,O4^f1AD+N9Y?T=/TC<<^R=Y3a-#.CE7Q[75O]96f,8YA[QdF,GX<(I#28DZA@.
CK1==Tbec2CA=@=/F9e3?5<&0WZ^9?F6F^@^I?^584X)eKf;J,VWgF42\^?JF,PF
#N70P=.N,Sf;K]Z6d?>C=_3?A_4=\/7_9]^W0,90U5^9\M:2A8XcMJ0SO6>3W=Y.
DRSXFI(\f@#7b.b9e8GU@J/\BPdOKObScfG#TBeX((>G?HGX>_g_abF,RLWgL8E4
2HK&9\0SRRJL+#O]B9RDC>13d]efVWZLU)MeI;(@44A-DO(K4b96/#./LbIVJZO=
??f+(+#0=IVe_=F\Nd+QH)]dOg1a0W?g:F6IdWQ\Y2E.T/=<45DBaO>fH#,+f-(K
X^WLNP[<E-9/OaN5:W&QQ^Wg=Ze3XZ/NO6DfCR&)J-TBI.?#M6K6Za-?(AGSA[Dd
C<WMYe6ISg\UGgMQ@A)U=bQ&?H10_aGUV_/eRc<U77dJbX8dSWQ<9TdDD0__NS@,
EXICZ]VK;gF6M;AQ7g1?O(\8Ge<ADc3I?<\65MRJ;R;(HD[2.V\EKdU]5^J+&6>V
T[NXa&ZVF>8[KE>LcS02\J7S+6\Z#WgNe,62QD:?\)&aaAfP75JbAK+TSMgU\+D+
Z>=#9)(]Y0X6:.Ef^WKM5cOC3#\+ZR(&_N?KRLV1+gPID:#K)G+40PWO9HW86=?A
6?_QGU+9V3BKb0;SIE.?A1)),ZSAL=F9SSMJaL3?SX8;>^?MQEWLD1(,](KfPFP8
B?EKPaELRRVLTO#bgX<<5ABU:9<MUW6(b.FbIYK1PX-\RJ?(Bf)&Y939+;VJK>:&
35JF13G^9#_c)ac9aP#>24SZZ)HO+#SG0a.Y8N:XMA8d4e[bU_NK7SU.f&MHSUcC
\9=AV+&=M=S5SXReDKF=D2Fab_,]Veg,8P&BXfF&8?MY0gF9:bSNR\>M^;])>27K
#?\N14dKJT&6UAB[<DA,B/3(@J9:B]LbDdfbSd6W>K(J]^JO(\EP[9LP-^O@A4ed
J1D,MGRNNdf_EW,cQ5+SbQO,EXP]P,Q-I?M@TQAG,+3\dG#8L8a@TC#DcA/>,2S7
<[#4E/0PX]04FY(=RCS:S&Ub1#c:1A/=L4T;.EO&>1d=T72G).-)JdA=JKO#V.<-
C5&@P]SJGV2;DHTP)Y?50Bd8]<DTbPgX=g]6GP)R942?(-[)TP/</EPS?.\3@9MF
CF@7CF^T>W4UXd7ZYQI]g4BZ#GE<(T7bGdAIE?1?,N^G;bQ@WZ0aPW3.,9OS?dQ3
ML+9EJaGB;bZ?=UPdWL_0ZPS;?H(C(Na\QCffeF+A&(TI]OEZ9C9aARGf4g=KDQ[
HF=(LB>e)__?T\B5CZ&b1,U<RGW01d5-ER?T>/>>E-W@;Z6@>F?0VbDgcYW0.7DD
C4U([Sa,7346Y)/8gMQL;FR=e1Ce-<WJPE^MbdUH+R\O5KPO77SJG-/@G#Uga[90
[A,V5XS2cV<Wf5O-PLKF8CMUC[Nd0_/RPAWA390CcP-X+2f0VLdDWbJEfN(YW054
[QQ]8_X0].N0)#Y)[FV\[L]BW<Z_,?[A9d-_B2V^?KaRBU@<eV2<J729d+=@[a.;
Q[4R(fN#d95J@QAf7L=aDf;(T78IQ_N)dVY.[V2,=MZ]-4&U_cc^f4+e>X]C,P#d
,7?H5BG7^@11_C+19dN=U-8XTEVB<NB/&1;JYbaZZSd0[(^@Q<;4Tf^:MW8GRf(4
RK>0WDF(?b4^Vf?MQ(MS6#VYfbDXOC,Ke<AXeY7WYF]/0W;GI]^e#(6K8:^84_S/
))9Y8M6T=3gD<F/6U<dU#:X7THW+g&C?@1NJZUK)gd3gD66R3c&)T2c6Q>0_,S+g
7G4+Q?e5fZ=[NQ6(W,4J);9^62@5d^--g0&[J&g1RdV]HXON[T?,CX8OT3fS3O7c
1R<aTS1+1<,X/1Cc[e_R85K#:,a=CWL5,A]&ARB\PUMgKg>Z6R=_2=b^Y&^50fZ[
K--83e,,4[/;9]MQ6D9R?f7_G<23CS&AABf8,#EJAG=@JYL2]F<,1g[F5947Kea2
+]PKIAN8:[E5f^P_>e#>5F]-g.>4V:cF+7a,Y-E4=>-dSbX4.6c/06DIVK+Q_PI,
-f/0Cd7:SUT)NPg@WWOH^?:Y+6@/L6fg2.7NPE2g(W#6f?5f5E-Af9^]B^_d-ab1
AJG&=b]S?LTWBZ4E,V6PG^[be<Ga]RI.IWZQSEF@:-]G0\TH=JP(7b@D_6c#(9/@
AXaOG(\H+/+dN,018_Q3Q5_g_^bG:D59XeE[AT:CRRMV.3GFG=W((>/BLSXHc\<>
@QEAeGcZeRWU,MI@P5IYZL)e9f<+VW493IH8#\-XO=6Q.,\+X?JT\NW?AVYA-O8;
_+E&+/2:TDbZ1\e/]d6E(.f;g=<:;(@ZHFA&L=P&(?8F5Gf7K[TaMG)7OY2=XQXD
.d;deU)^_;;LZEH>Fe6Y,;;D,&>d>a9YUZ=^UW5^^M+Q6G,#@?b3OXE8(YG=K=?)
+e42,S0f=JcU6OJ^G=ZgR=4AU(LU/M[N;69e4-b86A\D)CPQ_K6S9SV?0(5e5g8C
(VA#<U@NUBL/]8be+UXF@IWHEaMg1@?Cd8H3[/83J)^NcV^/Ic/c3dX1EKO\Zc[V
gG?>]0[:&.EIY]Y_RZ3#EV^0\<Ab@;+VF(NJ(MSYc1(^)&8W>eN3IOFRdSP]CHW]
E@#AE(N-;#>Y+6/0:+T5QO?ddPO:>DC<9U@8QLK+=/@=4g?343e10&Ad23@C(#V(
dOVdJ9/5&AYN#+Jc^>2KT1;,(5,#P/@g[ZN7UG8O;:7PO&?EKZ:e.2,E:=c6VL)T
K71O6S83f-3e6+6P\W\RWT>3>gH&EP^Q?MZcG9TgOR^0FF-I]C]EK[O_2>M@Z7WU
5R30(WeZ>Y.7MG4ebaQD4O6cY7eKdO&+S[DPZ#BEJcfD:1NSCgAK7,FF21G#0(YN
Y(4IWUSG=:?4N9G@e4O>9V1J#:L0W,3U)+Z7/@D:RT0]JKf:G/:7?MB^O#G/eBBL
[T3#98fM3(&[[7__=&6EFYS9K2.>9ae<U9]HBSMG?0>ZWW=_,84<WH>:R#)E@=-\
KBF#?9g]Z;<Id/#F1JJg--fK@0:9b\:76\+W5XON.TE=2:XC3C\G5^SMg1Cf1/7X
KQgGHF@1<+E;>LOXNV0T8(/5()EQ\>7JbZAASGB<bS>M]J=<gPA=-Q=G>+^CVJUQ
?fcE+8_\\+G.?e:X&>[gcCH_fZ0(ET6b&9WX&>RACGM&3T]-H.+[F+JCc:09A)J0
-@R+W[>Y^:4<9H?UcU]#96IA?)+US-EGd678f,SJ1b\)\//\6:#<:-@-5Q\:[B)L
7HL,1IG,Ve2+XW16J:-7D:=Qg>0(]g(Z3?[P:/PC:_&,)ZYB;^#_BB6H/20@>e-@
eENV&H7WMPbAYOP&RD\g(^PG;I=[\HVgfBN8Z-\DQ-MH1P&;?W./.P2CCDgMG:)T
23Q.G6+[;3NPB5>e2]X2.?G,4YYMe)1&A=J@9f_#[52J11.8^\FGb@?c]J#ag6R_
(M@LFN8K&bC2T1IG3G+P^CFFA=dOJ[QUX\b3&eWU<SJC?FdeWbX5Vc)JM(C?=BaH
6a_K:N-16F)SGeWGR-IM_U\0(Z2=35bVSF11B8T?P,F,cN>N9MCLb)NM.e:\FX<0
1XB^,6=Kf_ZTW>P7NdCSQ+GZ<=f8U&MfIX0[\85?=D^AG4FHRbeP:Nd/G1V][Z+G
V50#XHO5&5HLD?Y]?Ca/f(VDI&IF1bY;^8E@g4_bDP_DDLU]NYK7//<Wg^;Q2-R]
3.<5@^73KFG0RO(/MOFCHA,dO>:3PFZ&g>F(D&IC1O+(OHD<^8LU4J=&L\2,d^2,
R#V\XU+=\>Q0;=C<#OD;5#MAH[S1ZTC</9_HFJ(LA/S\(BG\].;L-.C>cRYG4?cX
R;W6L:>9fI+333A<4_Meg/J\[5JYNSUS6<IJ>\11aQ4[Y#.Z6I66Z^^&XZA_JC.C
N2XXCa0b;R^7f?378dOO31ZBgPYOa.QJ\3eb+I>9LPAPPZR[=DP/KKU,]\T<?eY(
1ABFF.UFY^WD.A<1e<D64\T4&Q3B@@U@;TT-]B4:NRFaaAU_47H[2\Q0MfTC26NS
U1bZYKI)C=/SR(9F+<.Lb:>E<\ID78.3&^MEACd^N2cCXRC/O^9JMLc^J?++MSD6
-(5<.SJdC_D&0+F_RA==MET3.NcZ)9B^_g13W?;^?IaVdRZ.TC&G<](6-cSb0bS]
J4]];[6?-L&^UPe8WaXJAL]8X\aP+4cU1)^]/?&(<_-&a#,@-<R+1_-\6DRaICQ@
N0YEMf1H)0RTIJc#.#/CPg-9F1#9CY6PA_V&P4f##BO.bI&5FM(E<3bB+.O1@=[]
O-ON=Z,Wa&,Se[YfX:CWf&JGQ0;=fWI#[6cd-A&7YdUQ=A/OgM3(\bSH?.c(;?]A
-0g[79c,@FP4cE:SdW1Z8a7g:+EF_::(J/X7>Lb_\(Q/[J0S[:/M?_##cd#=VO&V
+2ET+[OIf;0.d>3H;WE2BBB>_Y>[?dSga?Y^\U3,4C8U/cY++6:Z)I,6MT+(O4@>
NFc]GfXOLUX)D:Jc.(N0?8,R/4PT4(J_]WI():0I7#OXaGE>WA5?V<ZL>CTaPg,9
6RAXa-abLSd\IV4/K1H>;N1I@39T/SOCgaQ<#S(@M2FTaEK0^e]J55AA+V]C:eUd
aY#)IIW-g17#7(g<#bJXM[[PWNg814BFSNVV:T;P\G?>2aB&6=:>M5HR5+BTZ.5d
Q1R4F;-J/O?(W&>Z^&=FWMEQUM,SE50Mcc\Zd;NN@8DaSRQ/ZPSK3^3&8WH]>N-8
?GaCe\LU<F/RAfO]P2&c.L2)3Cf66C5VB<7^]DFM\YDSWfb70(:L1d&?G<c1TM]5
[d-e;bbU2LO@:3@0SfCgO=P5f)U@,L(AFH\XW5/g1DaZ6e6>@BdCI>51>J=H+<6P
McW/YCDGga38/MK/1g6RB4W=E6GB#E8cPg8?5M;4KT@_g_+<\D>;V(JDTQgN[^7Z
YVSK=W4ND#BU\-U;EJ]M3[,42I.7;3_SVV@F;A6W5]Xg1KE[<ME)\JF;=egTY?+R
J#3O[YZBO#.7\YeL[2Ca>7:HYeLe,WP#CE^1dH)M8(C_+>UYBVe86AK7b?3DEEC+
-8U\/QbbO><E@AUV6,+L;Q(,\XZ.2NFR-W6OH0CdB^4FYMG:A6F?>]\\RORFWYWa
+DVNE]KOeO>CQ))_::W;.DWV5UP46.S,ML@fTL;agYJJ40FA1-;T7HaY_b,d8<;N
)H;C,;cMfSA:>gDFPL<W\4D@eB&D?&<b>=3,[1>RKF](QT(7Id7H^ebeFd=+a2dg
J0+:5eF@<+D_D(_?S@03FFY37ZA-#2D+U/=1ES\(?>H]a?DUdP:KH1\_[#)NLJdc
?L8#.d&6f]HKQ<^N\.W8PAb>+^ADC+ab82L/0VV6Z2OAg&MKaAUEN9GL)S0750Sb
3/U>-MaaIQ^XA:>)UG9=9.Ia^DCV\]./X8;d(3F/I9-1B50UDWW)6&=Y5b5KMB9G
]fLBH6&L156]J/NAe;#(F8[N;M8>YGfZO/N]YG&0_0UNeRfKJ5@9A/=Ydc^XfEcF
;ZYOeTd\54E&@4QGG#7B:52D+@TdSI34#GF\LRXS?@fe]=<M&8]\7TV63S&V2O:)
L=BLV@S^BF?O>VZ_R/E4fG,KM_52J7SS)gEe)8SIT,?[&9U;Wc3U<(53f6/26^00
?HUD,-L4:=4-DP4J/J_N@eBI8;d9Y/UJ3&JEB_HdKU6MAcc@8eHg:LaY_E\WQeb#
c=<79809&-MUD97A?gKHXE3)M.@e(L?:&deI1Z#]3\H#E>]Vg[A]-Y=Dg4B-8P44
&/P@Q.>A^-GY>4[ML6c?NHI04^T34#_Z=[+^(Z<AH[-M)1?Z?QWP?Q@1DRCOS^=Q
^C-1a3C2.?Z[4;6;@H8b+Z.KB=L:T@7eEGXa-/^>2;^RL[cJcDgRK;>@47C1HHEP
D/V19eOMAW<#g<\-a=X[.)3\(c+^c675gN9A&K+JVYRIe44J:TXZeJE_)PZ6P=&e
IIYaJ2a369#DD=7Q)QdA,P2CJBf?[X<:6(JA)^I[<,Q3S3,4;>[#\a/1?L_.;^:O
K^0cB6>?ZYT\J]-FQ2847?4?^];#I=g5/]#YSb;EU&e.L6&YVdC;O8[6f#&gX@.?
E@;[Kceb.2GM_JXQ2((3P991aOZY)#4d&>]RY=21b9/7cg>?=_&KK;:D5+.BLHdV
EYQSO]Q[[8GM;:.g8g<:6SH)QYFYLLTU8fW.<0RW3+gY)(J>W7(+.K\ORT>#^[.c
8:YP\GLYV8)6f<PeZ(c)GgG[)0@87=E9[9SQ54:C0X8cZb#gL<Q:&O(dIK15Qd+I
T\4ZP#Qc0e8J8CUN_^JNa50O4-V8=WB?[IA3.6<V^:C+0E3^(XT4B>c/SH6cR[++
W;SY3^cX+I\:>g<CeTBgg7IBEME5YTBdGY?aNJIKGVE\=:W@,XU0Ag=2^g[M@1>T
[,0(Sd]S,(;LN,/XVP>M/e(R=GCAK,\LJPZPEg+M(+=#&gA,VZX3;#f>5M0;R3,g
Ab^@]L6WRT(CeK.U-/d;K9DUbHbRWL.9T7ePS<SQITL=ER,?8e_);PIbO[XG-TV/
VQ9cJN:f0,I.X:;aWUYP[.M186+V(+,TX60f66(I3c#;W03;Y(\5E#1#,MSV\H&<
A@ZWQPg,A;<^Aa&aTJ]df:@1>A<cA#F8/8>EU^2OX129Z]-(>H324C62?(ZeH=I.
_(?I5NC(F+A#f1(H+6]+>d.&DC\I#M007HU,S#5?4Jd[XPW^Dg=MgGLI\8U-b(&/
4aV5@)=AQ&NL_V2:0.?fUV8M#/W#J],(_?)CNRS)TdUg]KI0T6^53+L,;;MTP&?D
?^0&GM7.L_KR5E5[11G<Z/LLLcV;eDb\a-(#2=?DTU8,KJ_7T@F=cPGG5]]B9_B_
a6O<ID22V<[<X6)][KM,58Q9aTXQBQY1)fP&<BDEU8#7&(4Ug=g4>,YT854[N[e3
CfI)CLKT]HI<:EUX=e_U0RaVDg89Yc.SQJKf/[064PADYC(&CAQdZ:eNY>1K:O6:
cPc0A+(eJYDUL.A?3L[D@?CWOD5A7D28eU_J>,EP=:0;+U+69>aeC.[03OA3PZKb
S:fX)_B?TIQJ=Q0LX<,W+H3c?V8.Ae.Y.P[TWa]fFB.Sb:cG/ISg62D=N8@HY?8Z
?))=DBQMb2/RdZe3F/T-O4JU/9(OL_(X\0b<T<NP\VI8<O?T?5ZTgY?LYRS]10R&
^D@Z(=.MV4#SNS^LJV5#NG:3-Uea8(NOc0W/WXZ_L9_NBSa3025ZEc8[([,,:S)E
5;.,Q4g5Z?J_]Q1Q5K7.==?U:X=(?Z]SP[6;TF\L>]PFd6ZD<TV^SYFS@?V\;cW-
M#cd/d4#D[]VcbNbd?4:@2Df)V5fbIN2KXF3DM[X_9&VY&QAE\.b&,BJZ2@Q2XO+
_E14(831Ng_0b>1@)>TB^^I&VZV]0eIEB)=1,7I??7Igb)M)AHfOfPW\U<W\@:^E
bSbZ008FNF2829ec:/C?YQ<-,^YK?V,B9A4KPFJ0M00/T?eab1(Y+?>3T:Q<L>6c
d.N<[Z@AF=[eH?J;ecH_c@:-e)/7fY:W6?U4aG67fRZdLScM3W40B:M])C6g]@X&
dE;LcVKRX/2^Mf,5&TcPdF&_0+FB/P2[ADZ?OaXK)+G_48PA<a8Ng_LZT>=W)Mea
ObfFLf;BI-fI_5@>=\<S4O^_>7f;1W;B_72#NM>3QUOR0S\@0([X>KP=Z/0T2]2G
^233CfcK5&793([;</HgaP>,WF<UIQ;5SB/f][-XAcbETRaH6[Ga])#\ZB#7DAJV
<=@LS5N[EZ17cLX\#]Q@]YT;:-<6f?)N+2[gdVP);R&,>QJX9]L?-]QWEA#>g1L;
G]V>W?(9DP315KKZXD3HS>eE?&)d8eM114Xe5R^ERUJAWHX3Q,_)O7:<ZO+N?/eN
48>H,)4/_]eMHYZ,b48e^PB(3#H41^fe9ZI/B/V>I\JJ28JdX<-<H_]3a,.TI^9\
DJ5]>1JagBZZ1?ec2gH.>B[K-DZ90H9,)+K\MXAP-K7PKS>3))UKfZcNMY&a56Ld
>gB)K4I^f?Ag_cd2EN5&K^P_?0\C,JWSg<LDLN;VW+M^HDND,<WM(I8VKd,GP?CQ
;6bZ^3]1].>Q61<.PV-g6QRD@gKV8^)2#Bf+\6X]2fX20(4:):GI[b;d9Dg[3Ebd
\1cLL^4#K3:d<>c,T0:F\P<7GU1?1A5?U&DA^a?=6b&a+[UE&^b0<S=4H,^\\P;E
U/_adG()_=]Y]38TP3=NbW:5WEKOU.D=XJK87>:QA7C-Ab56>ZL:)UPe&dWD-B+]
LUD2L9#DOP7@;VHbV4.QaF:6#+D=7S/QUU54EFBf(B>?YS>>)Md<eRPNc5ZU>UK?
fI6Q/;IdV\bMVJ[e5B#>\425EM^g@#6<P),LY#WD7SQ+U?d[U(IUM@O3+C>TaX)g
8c#+PC68TO]N0)_M,Y=MR;S+^PU(?20bf,<2(92+/L@7_?@,(g@8K-,K.I.\\QRY
E7(eH15Oa/15>@K3BXgOa9M/K2G-\N>WZ)^abJRB,8Z@#[J;FDU^P1BT\10QEd0e
L/4edeIB\N3(DGYHLbG[3TL?S0&IUe8RSL4F9+O=,,W,I.4fIM<78dV83[T<0?]P
PM9Ff@&]Z/KCWU8ID3aM^<f9XUX8:T[>;e6B\RZXU26O:^C)TI,b5PTZ<NE:_K6M
BK(;&3Q4?AZ+4cAd?Q0(46Q@T4&YEGePG(+Y2X8GGA51RO8Q,HLbK<[d^^H6@H:P
=8]MfbYBNgbGIaM2JRT-A+g83Hed#.aW>(]1,6I1[VDd/(VIGE(Dg1>0<;XSY]X^
1,::PV#R:^NA_(F.UeO&eVcP?)#VR09;X[M)?H&9cC#f&)db=>;YZM;B]b65J5(U
R2Ka27T]1+D:0]Q[]/H\KHY;<^#Ic@R=;X9I(OFLJcAbF/(IA.[<]+0=IdS(NT]9
g]R4#Ib0\H+1;/A:L&A0Yef<.^-dE5a8(NaU,B.<5^RPb#?b2=R@OC6LcL\B+MZV
?P;DE.<ZPM@NO_5Tg@eZDCBN=2;&[5S2<>/2=BBXYD[9a^:[N[=J9C<L.=d;_dPe
N)+]83[D+RN(E-JD879C?8T]K4DQ+KZD>CPH,\d18NQZ0G?83fJ]X_5.2(dC-BYM
62d,ZHM,.;#B0=WV2,aACH\S5M@AR@TZD+E71MN]NQ]=DC7VAAZ.4cLcf/GB?^O<
:GE2@3T\GLCC42O?3@5b>[<d9JPBA+B8(ELfeOgBWBedgKFIB8d2@QDgcI)K>@YD
>-PC&R)\_QgKRNNWL66Jd6_4=>g+LX7S7fV5F[N9KV/NVeP<)D>3VT(7WT/5dB?R
&N7R#S@Gf6<NaMHgQA&,#1H+?3JG=SB=Xf@4ZO]B6N.S/Z4]b90K&PQ5L7A(40#W
53CW9e@e649QM9(JO4//TDV(;cK,,\;;B2dHMG&(NeT+,1WL9?.>^(\?QZ#(N<:I
AVe?EK=gSaJH3[V^2+:E@4dM+FBE.Oc.B:f]f98FB]QMLFW^Fd.Z.;aNK&+VK\Rf
Qd/)2a85,M=O(9Q320a\[Nb0g5BWT:C&KOK(\C()B/G\-YX.7Q[:,2LFG(0PS@Hg
X0O)e6TQVg=DdJaG4?De2JdEfYGdUI@38&E]B_dgG2BJgOUZ\c,@U:=Y-(5MB8^8
De?8bRI2,J^^^_#-e<f-Z@b)bdN,(LDc3O;2HL-Y72VMXfeX;YZJ\f=2FgNd-4[I
/^Q/19<::ZO&a=9YIIUQ(S[?\7.8;TO.Beg)6MH6<X#IfA.\X)-RM+SeA5@36ZVa
f1_]4cQW,a\[S:>8>f).-3=EJZ@8;I:2<fHRNd4)(X(C32=gN:b=KV8HKPK=:,@g
/ZCPBVX@fO[EENGX1;#63B]EZT#&CAd99_YV?218,c4>bEB?]>FL;;B2bUDcOM#R
SZ7^CSbG3R2^[1&FJ-cXP?>)5WN0:0<6e[@cK5^eN4-A]>JG\UdQcZX:0W:OA4XP
HC2)N7XC0B:4OAF^8bGXMA]e+NbP-JS9g_6H=0>-PVJ-);VUN\^XE5K&Ja_L-[LA
X#6+Z/MUAe]Z6_Y_Q)F.Sd8g-4#8c83PS);WDZ[<GKR2?[179a+fd,5.K0HJ_+\Z
5@V^CGSED8e;eH7)IU>L=WaDAL39MR/IKCP:[.O)JZLOV)g6XBd3LD)e;M77X7SI
V+,]H)H09W#W9W/206e@JCed4a]_=PBSU85TO\(6:W/(2IZL#+c)JPFWXgY^D>OS
a/M#Z8bG2]3V&?=>+&H6JRS@Q&IV439;)O68dgNJV9>>1U]^)gEaLM<fZ_J:6LI4
IDdKLT4(GRS0_GfNg<T](f.V5H@:-WE+9AAK3G/&JCg8>bJ77ObIe]E^g6O8f^X:
UZ5L.\d3P01H3@^[(ID9Q49K;T6IDS#?NLF2)LN:)(Gd-V;QNN/Y9C72Ea:6g,Y@
]-0FOf6f.C9UeO^NOAT2=_.8DgH6aV>fBM10\<5QOcGOf<#^S)3d+\3+@eUS@0.b
+3U]V/]<>#,HJ2\J7]22b&Ec^XD9<]TFf[(E5bCag8Q\G2cDJFHQNbEdd,7HDC9/
VY9G=N/I+_7[I?(,/+S+24P7>40-5F>Af,QLI)>5b5.W5MHZ<?I9L-c>WYd.G[GY
\VQ=0660EU<6853dLg#4&5=V(E@/S[77d_-:YLgQI=./gf5W5,)#7?3^\Ja<>](Q
N6:7O9_HP59;(,+-OBE0UR;AHb::(9IT<329-JIFJ23Yb#;T5X6Na33U>V)#Y8=1
P@P8g=/42CQcM#5H_9&]JaJ337[e@ZHQ+Y>JV<A[:)6GL709Rbaf#UcK?Dab@9=K
;J,F+883@//6GWDQTe4P5a?.^4WdK/e&>3.[PbdVbL8Cd,-Y(W_eZ9D2cUQAAHd8
]J4<]<UV.?d\]@[2>E7b2,YA6^3\CTZ\ONB>fPZ>/\264L:F;gQ7PS:FF5>bE3LQ
M&2T@3-/2(g5g(VQ[;C.)M^9;^]N>:fe4AB<La:FX(]d90[B8(3S1YRT-OQ5gYa_
([RG0_1gY5E8acZ0(T.(-&ND=Tae-^ZM#81L:NECT=JO@MZ&]1?fO)]8O1^RY0>^
7\^YbgVOS:??<f2N-Y4],F3/>Va1],e#eM@Q](,WB[LM\U[4.<W9daW;4&\D3f=O
,gcC)\I0.:d([e-^_I(2[\VC7&WBR+9bWRc;g#2>H4K@B9X2d)=,5Wb0(NIH@:/>
4E,C#K;AG2XM[>#)HWJA\=+MK.#1NFO:Dd1/F]SMYN=L\/_/T5IJ,>C+^Zc6Ka@:
+SXUHCF[E71WMXbEIKEC[&3)eS0(C_eCMbb-3L;D(^6P4:>:6I:11QL[_2c0L<7e
g<-SM:#CAA\^4Mg=(<d=^37FT[fM<Q^>ZN59#c#;A@>TDDOUOa4SA8B.5#KH_.^^
XN.FcIU:2QEO.+^XcT;2fY<cDX,(Y/XY_+?=HV;O??,C\04;<Q/V2.T_WRVHN84@
CGU)KAeG9.@<C9J_4]3=0=>C4ZOfdSN<&?S./E(IT.gAe<2\Z976A3^A+,G,]I0E
9D^6::e::8W#REda_WARGOSBT5R.DO?X-]0OT+^^/DJb(U:PCC+B36&1eW<F<ADK
1EPI8Hd6ZS4=]PU<6a#d/8OIf<g&]\GB,RK0>3)RP>ZD0SRUEc44]#XOTW:.OacN
N7/7==VTVV1-_N;f;OdH0O@-0fA]0]903C40E32UcGD?[F-6V6;12:#?,,4A.AfZ
X0GMEXd)FSSbI8H;?Gc[I937bS?#;K1IfNYY/^cRcK;9<HU#EGY?Bd_:66RWaQXd
:Z[KNc1=FR\ND/-N^[0gM8+_<D(IEbC(O<BeTGa:RdFS:H.&8,e<>F>Ye+(4(^K1
M?YKY]B&/M.WJ/cHVM.9@?=UA1K2(e3b<1b8VMAIENYCH_>XYMFMZEFYI0K@OE6&
X=S:R>f4RR9G(&ScCLC/7_TJ-<WeOIM+/2R-A@Qg93OG]_<W^O#_:UFQU6Z,=^.?
DBVS?OJ:&0f8)[0]aAcU_Tb1;gbN/XdGZB2g-NSe/MC\IX75KCM53>GU+e^)R-A.
N<U7D]Z>abE+0S8gC[O1M+7Q25^G;OXEA1I75U/a0=30a-aZZcc19Rc2)(08.b.g
NK)@W^BMJ^(-XG30E(cf)_+DWF\QFd+.LYLO[MgDVHP/(.UeUa:N.HWWFg##gSf(
Me2S2.G0XTHE2-NWW7X#:VMLYg?=BaY\P-V^f=W[+WJR=RE,+5-I3QUV<PZY9V17
4Y29^FE+(;,b70G)X<:-</\EeF4[dFJR/@_,#66b84E-5G58^X\ZGK3338f0E1<O
WdZ_RH.1;[@DQb]I\MRQ2HCZZQ^UFP<T;W6/QQ.7-Gb3e,KA^)@YAXga/@-ZYH+(
f8gXOY@&Fd_RP+eZG;/f<c:P&a^P14]L/,MS5Y]PUdc/08.bdXd8AVL?<B1)XTWd
bKa<+cMI-:c#9U13,FJJC#,:]9.WC\0OeU#BEXNEFb+L<O6f/Y)-cO<>+BQA8+43
Y2>2/)A>]Ie&3-<N,GL3N^_eTY0d^FFYcI+]Ba#X\9Q-RYaB?_[S3Ra7>1Yd>c;-
UId;,9PaSBU.)3[\VM7b2/[FNg;@W];9++,JAeX8UW/)9TG>KI/V1+>ENM4/cB/,
>0?U^0V2MK;&-R&WB#-,R?6Ff3SGQS<.e>XEgbEAYZ_@IKNFI;fGYR6RP^+I8cQ.
?f45bVY+g,VJ[=PIXU?QTb&RfFR#XPJ#/+OSK-RFGV&BG_bC;R9B+25F#CIOV5MP
3J.LU&L.-9CEAL-f9EVMb:SUSKS-;XXe4OKOP#]<RD44]^D-?;;O\E9,G0^>C4]3
=(?BCXNDObUY]UY,=5#R55CfI9f/OeOX.c59<>3U[bb.:Z-=cfXNa5<D;3ALD9g<
<QD.,07/E_K-WQ7>9aAX+&7eB7\(\76cY&][>g81L^@4GdSg2d)IWT1OAXceJ2D)
&V;LWBe,8L<WR?=g9R_0d(2W2J;5b2[8H@g76<14]?O7Ka:bZ#CM=3b7-)K<Z/K[
48PO3#[V8KaP>V\_#b9H,\,IAKX+P7<[]<g)FQQYBT>Q)I83WfY_fKcH5Y-Z&b1]
,A5V&J1D0eH@F_IBOM&K+Z&47\,(b48cf,;ab25,U38d)3G(B2CS0BB&&C4<QXXS
G-\/G,+;XI(+(Fga\OVeJB=RdJM./:GLdE^C2(NSL#>=?NR6^9[H<573CIH(+^QN
,0cU@X\-<N,KU42R:EYNC&+66;59MaOgG>U^DgW;c6V.NW0D(cP77<C+]EUV.gQK
b=4/YUgAe9W/Q;JP=Z:HDcfH(<?_PEKY_WUO-:_cQ0O44<(EQA])M,G<9WG>@.D,
2f>c0?NL/&QSHP)2D46D7&\,3U9FNF(MEY:<8O43e=1LFd4LW?GP>U]]2E]\04R^
C?7bXO7_6RG>\Y;\9_JREbVF#+7QfKW1eGg[@<(>+32OG]OLD27SGQV;/AIIA.-]
\+2?a>dR-]fZ_)GE0P]96c1OOYS90Za:+@\OC7JDP]C2ONP<V9T@E1,bH\G/X59P
abQ//adZ_:\HX_Z/G?Gf)VL7@_+G,O&W3<b&^YJ0S(,/eN.agU<.X67PN,<&F7f&
>IaBcZ/+#/bZ2=O5CWJX5O08CF6POJdC=f\IgZC4F/7((]9>IOMNX@)>c.58cV/5
K>?)])I>SFV^87EV/3\&_M;:1(X<X-B^ZZSZM,QS-OReADIWBI6NU]@02QKWO&)5
R)8E)b.a1E20##Pc[d0C]C7AQZQN_4K[Sa39O@bcA-U[ACUZ7?Db<.A)P56fQBde
7+-TM>>EA#J33TP>eb@a3d2)E(,Zg\RF1bc1WL)Z+ML6\\7[9aY>EKbC\N[6UNG#
O^5W^:c9D&66YH:-D>dZA:/.ID+2YA0ZZCO+[DX3-G4C^EfF:/bR+F9K1bg\N.NF
#47eC_>1-9I;P^(BR:31WY,OQ8J)S+(,K^\5FfT5YS7SG(SYE-/GV9Z(;cZa,cD[
[Bf&Q4\U9]BD&\0#@B5c-\J9W,+6D2(6U9Z1/5#[82d7NZPd\+?4L91WHWN2A64?
]Og;Ac;E-9a.#&,9J-&-f@KTD0EWOE\C#Jdf58BJ-fJ,2)FAV,R?5=5]YgBU)]LH
<^Vb&D-?^PPY/Q#Q?7,<@60#6@V4gG/7\Vg4T22-d<+9a[MIgBS2ESd0\>Y8CNU7
./3)\[T5>Tg8L\c5VI/bVN3ac8,#&JTU7b[G8BV_Bc6@R]WJNR_?geG.>@EV_KbC
_E=dQfaIVT07X(C]97(c(.^8II(Z/WcAA&2EbV=L4PSV/]?R1-&=IZ6UeA:I.N6?
PE3M9Q3>6Xb^EC;M8NE82>gU3V0S1N7T^FOA0O+5>.+>3#T8X+\.[/;</]<[[ffB
(BQ_#5f9;E0+bcLbEgfg7NYA3<@+.70RVI<?&62bF90LAMa\+CZ(IM=)&Q#(LM9O
W4?fV,9L6/:&9>eMQN.U,C&+0>1,E(+F)O.OH_;eP,E<&MNM?J&3.4Q&D6J/>>@Y
E,V]XN@FC8HB7#d1^:#FdL>J(84IP+aI&R-6M?,OC?)DEQ_(CM4V>aQ4OT>OHF;F
=f#KF.5E2K_>Kd.C44DV)b:_W#,C-)fPaHPR_>=+NYQ:.#MVO)4N2#NTR4#-HTYf
MOZC2_bJ9#\U:<VFA:;SY,CKXbIU>YHgb:JFWBGG/H20.3@HR5^eZI3R.GaWM+@_
?0JGd/W;?Fc4/4ESB(PRg>JdD=C>2]>aIMb2.:>,_(3>^]R_Ib<[H=Q=^5C5K)/8
OIN#BL\(2M&UE-1V7_2UB@S^[/]G]@2HVY?b>4.UaVJ)\ffU(2^fYM\0G@)a1O80
a1P;>>I5X3#D?ZQ:ZR^NPdcQF6WJbRY(J:8_99]#FHL.g;?g-RM(RHBa+e+._T)b
XQ/\bJeOA5:R)@,WR.?a+0I49;e-(;+f9,9K6P+80X/2OK(F-AM]8XW,B-8UddLF
8E&W3H?^<GWcfW/-&d4Ab92YB,3PZ.DTZ;@gGe>K3S<C6SQ:c=_H;cd>9d2R:45X
&+MIZM<4E>93)-8FG0[6WM#W>&X:2ZO.2b&<::Z(C][D:7H<GB<Nb-:,EL6K4)Ka
6(OFfI\g#-\ZNLI8JUL^_2P+A6J=X4-XS2&TV[-A7>BIS^WM+8V@#50R/^GPUP]5
54aeV\<CBM>J9e&<,JLM5>.0L52GO>L6fTU8-^OZ9X6\HbJ46YP2c8D@-b0(N5#d
]bZXfGT88_3AfP.D1a-\ELVHAFf(_PdDN?^8(IALRCCfRF3gZZWOEU-<FMWQP;f-
^/U\Pe6bfW>VWYQ:)dAcAZ/(,a,#>/,+FGT>7[>0+]Z=5[817FM&#1H\(YM&I^_S
\:5[T2+4ZR:-1J2;)FfB+;DU.>Je#8H[\aM[K-L>86:AU4eRd0N9^T00CU.=PXO\
JdJAK17HXJe#eMO&bS#69RNMEP]b?-/IOJ_,.56[\9#&Z.=8X-0]Y/gS9H0TgBZT
?AdJRb+EY,;f[2fY&c,+KgEW_WVCN?U@GKgIJOGd[(V,4A,<TTE90T+?+(0d7+89
Z,U5&AR-.:fEHEON5J+1b@9@Z#>aYRbc68J4c9Tgg>/fH54O6L>E8K:Wa&8LQ0=X
^MD_>\,QQ]eL?OZ6^?T&IDLg8[=:dQIfF(+CLe_^cQV9C<(Z?^SS/K3fa].LK\NL
?4R>66Wb:L#Qb^VYAAL)SVU:D^P)(Y=G?;C#;-(N=d<+F91/>g8:BRZRXdbWC,&#
[7YB/:>^VN/AK>8f.a)VJEI7Mb:T-.U7Re4JL&+T>5?Jc\37)c]IFa<E(#A^^0P8
AF0([<(295WL]7<FS@]IRS3^+C=A.\BD;?2>]US=&[S844bga>WeTW:cE#U6?G4R
b[V-6&DbS7(fF\Sg&XO5_2IZ2QPLCANPI5K#H/\C?TT/4S@0-@T#]7HH3BbL1X,E
E^WVT]\7AEGO3S&g+a+?OM]R]-79&LEe&M>+CP<6:20R?a-SLA<U=]f3:<A8=D(3
d-OF]V<N@dBK=fTP6-E.FUX@6T?:1RDL9JCY>LE\28FX)_U]7B#+8:>9TRFC+O>+
P3D?a3S./NgfV?&RIH,g37L]>F;.cdX>YfH(6-.DK,FF1/)6Ee6D2BM@GB(HO<S]
e0P\^&X41>^MTICbFEe\Y2Ne6e^Y_2Kc??GES-/F:>.AAPWU1C[IO+/6(?]_I[(d
(a8Y?9/a(X;TK(dXF(GX6T;#)]>Ub,[9,V\-;55-@8f6C-BFR.GM7N9Og9N0(008
aa@AR2D7Y5]583Q:gYOa<7O@UNSc>A-7EH_CW]C?0c#LDD9CA_]ZE59<M_TJ)5LD
B&O6-&Y6PfR&2,Eba\2_HD,7U,,I7D=<ed(CW@+2gB:bCKP.-BV-WE\;<Q]IOBO)
EWV#XU<IgM=ML)g;D:AR7]T(??OXA/3abTC2N_P:2f#cEL:b&T4f2(LcIUd2AVI_
A_cYgG\]2BY6gJ)3/Q:#J_SRU&.S/T.SLTLCe[6SJ:JYZG7XgI_:^cdT6INZ1T[+
H5Q</,(_A:.Dg[.eJQO,QTDL2+Y)0>g5IbP\FMY7).PUGZ-Ic]I(TV4TC]X^8IZZ
5K<>S]GTRRcPY2WKfBM3WEM(=PW3.=>,cH0?K4KZN&UaXL5X#I9@WLOOENUP.b]8
c0-)]CH_1Q+&;;XceZZ),BaA@\#GU#C<;YJ^[;+d09LM30f9aP\27MgO>d\24ABD
PN</7)Gb<P,\gJ]WN)>I[.LbNT.^9fO.K[7LfEJ3SE<KHf+J-5JRE?[D0G[NJe=f
TZ?94RVKN,G8\ASXb)&fW>[H4-590aOec<=eXW9K3\3=C[)0A@N1_N:PLN^&O99:
&\\C7<\ON+Gg5H5M/UU7,)IX_MKC[_c=4c)EAFeITX&(_DR1ZK:U9OU[#K<I/O+N
gJ_5YaJCg86W;K<PAe1-)a?P5-RdRP4N1TE;gJd>+f>++&0GMUTR5aT]@GAS;YcP
O;O^\6P5&_T#OF>Z93^/-2R3fZC.0IfR[fZ8@[\T_@g@c>=]R3QE+ARF_=C3R1T[
5-[<=Q3URVVX3B8T5b)ZRfaNaCcCE^-X(?eW8>P+Fb7E>>:_(Z-0?VP11Y0NJ/@>
-H/^1Q5A/?>=_b7R/^L\7/O#Ce:3e:/:e50F4-#HR2CJbTc_e[B(YK\#;aV>.1Jc
[Tb7.:<1dMb[cJ6D(<g81_U=:Y[[P44T3dQg]4Bf<DH,[VH0UA<e9d,XQaN;/@_P
cedJc-/657]\Ea(Y(ZS-E6@;E)CIRVF+9RT<[COVc)__/aTT[;d#R5gHE52,2N42
1.8O;^N2RFWF4O+2BUB2)BTg&cX[ePU3L+I(d0E?B(\)(^TfdR_WJE7-YZXY)QMX
W:d6QMGfA.NX[_TKC_)aC]](=[W-JUO1R;R?19Pg&DE9McUQ/:\X]7)>HQPQ\_N.
X+b>4JF#4:F(OM57K>Z+,R4&,#<eKG:T3^<&P0WFX?H:[&HWTD?Y>BPbA<P-;^[X
BJT1d)WfFb::GME[C]&8e1\N+Q:P)XXB=MaLE.JA8-_E?TbFQ2/ZaXGQT?J#-OF-
>]KWT(U5P[P_G>A06@+4beQ=X09dFXAaaN[B1PTASE0OT;gRU9#&GJa)A;<_\UFf
35Q7>2<0g7f/V#^@ZF:V=;<PUENL_IWa,.,R--R@7d5aCQgUUU8VRDUK/5FJN\d6
^?6ZHH/U5L1TLfcAJc:1a_K<.MeWD)e<\,+&.HK-SK7TKeL]@1dB2faSIO>R^&?S
T+WA@H+JNM(HJZ^D]4V.A7/>O#KRT><8-W9bY^G9D=C<+K^C@B4=ORTbD\B=#?Ja
84A,eF_4NG-6Debe8;GfR7O4)M\a)J4SP_8J+CNS_SKTDZ8U0;IFN8-1U-Lg1IW#
J?L)eGZV?IVHN+ee59&<F5)8QVA35U,U&4I/#?Z6ZVcI67\M.V_EL2fP&:=?\/]2
ZFSHfDNS5@HDZW(/_GKdP4W/Z91TA__@5/g]D>BXM_g)<A_U^5C#N+O)H:f6\M7d
K.-IPZba^2,.J6@9M&P:<SW-:8N5Je=Ca;6Z<BPZ2():UZ__IW.8QTO)DJC&)[U-
+[?CEFF-18?NM<Q5UGUbA-2L7<O3Q&QIH>d:F)Xf,;9@;IR@(88c6)3SbQA\9WM#
??6[e:3@Y9RO;S/5bN5//^SdD6:AAM#A@Y;@C9eLUWNNM09:Rgf:QY\,-5\Cf53e
eH3_ZX0SS2?=GCS^O=e+RS(I(,PZ>3\AP>#SJIXb^_#b\CWTIdHDEQ6>.5#b[C;g
0(PN.e[NC&caNc#Ta<RA;35UN[&6PW(a6B?-(.D^C0.793TN^P1ff2/KF57bDD@+
;2XR)E,a8-R:eXB#;HYRLf@cX#_e:,:=O:_4Qc+)Q,^,]YDgPN12J?SJZ+&G3Fag
==/<(bR[KbAU,1KPONC_TFN/Z?J2;H^1NTD-V(9Tg()2S,92dS.6dQ?+1+VVSdZF
ccfdf=S\D@-ZTLU6LUX\OdJJ6W50F8a78)KJ1\84/dP2YT03S.@=.HC+aa_3XC<N
92[U>]YUff](VCWM[1IM(-4M8O\2OCH#FF1G/S/67KAY9.SLe,=@55ZIKT;e\Y?#
8e6^#J,M)6LT3_b[(cag7X^>@AWeg[\RX[VaS6e#d&6Aa>L<IH,gSA3b2g0O]4\Y
IR+(E]?SKe,f>V<4CN)@EUJ8C-;\Z;#)IT<KC:b,Q_G1?WVbKJ+,d>V]C/,\a\>G
cOU;1TLY6,dVg7E)MZW)8[4JG6J[G#a[3(6gNUHaOS-Q?:D#6.+G1R\-AO=e-<78
\P><YK4:VNb]\G#I)3<8-_)e^46OMC0b-1YS8C0R_9LfN0aP00,3d^[B/Uf6=PFD
/\f07Q-)#I:\2C^W\I),]c]T6]=.6cE8.B&Lg1WXCA/6T_S/#c;]d5OPQCTf+PPK
?8KP>b@3AEAQHGdW^gQ(LN^CE&3[dI+XL?H[NQ6ML;0BFJW8,D)>,f/VaRfd4Pf\
(0+3\J#f>5J:&/6-3=ff](GfGCX8,@U-\H/6&g_fN#8fX8_K]5ER8HbWICY>>Yg7
9bEEOXN1PP/YEA@#/SKA@\U4,eCO8]_G_D8O9dEOI8RZ]PVMGM3SS+Of)L:Y<]/T
gZZ@3VfZ^/e40D[PSQRQ0-e;MTF;Z@[C9,1>fT/a_?&)4)OZVeZfOPZNA2Bd/DVM
EH07.:P@b-]7I]/\\L>JSNAM=I6JDR\?_eT=.4B;\-+0CK=GC?6POIIYH4,Xd_+3
e,6Ie0WBGW:&0695BM?I)DPH/]M5E5SN&aYAGP1V2594#P.,c30CUSb<KHMfbBEg
:#4OE4\4b<gTTRgDb?#>[4eY6<M=)-_+N:MdI&OO>H\F#V7e,+:a=O29,Bd0?B]1
6MC&TGF6^ZR9,O/6@a;[@c?<4?DIQH&<-GU,Vb@8U6a=-?gW.+fX97)0Fb,b(C5Y
S0E]g/_)]?.=>_VHaH@5OC,1?W5,,7M(-.]QGHVQYF?Ac2Ldg2+V:[,JK1P_e\eP
+K=;?Y\.7G@dIK]0S<M:)#9[g;2W[J3EEcKBfD.OC5=W?O+fSgVL-0&&C9G.MAG,
CXJLI0_c?:MN?FSI(C\\QQS0,f]\gFe>BM,GQ.)NLYbQ/CBNLJEYQ2#.0RBE8T1N
(E@dP4YW9S5;d_IZ:X.(=]]RALCB9?M]\ON^SfARaK/.Q@4Hf>#93TU.X:d-X9Lc
Z;P4TT;cE]_6J95>aLdZTK01C8#JgWOU+YU9N,0VKKg^>DX;56UP[@I->[OX0\KB
JXRV)J2GXId(IA/LRY>R5):GK<O0#&Y8>1WKae?+@&M&Ka42)0d[RMST[HcIX\d0
<[F[#4T0FN-gJ/1GE.Fe(]2M=Y83TeLEGP1Q-05IF=)U@P.@ac(DHKTT4e\[]W=C
cRW>T[B&C))M;4LEcbXd2UQEGI][X=(?Ig:9-SN1:&>gO?#+^=422]\5bF#MX?.=
>9eSE49a/:C#DI5E)HY5&,ALMJL7LN(XaQ7/b/bS?&EF/c>52):7_B]c;0@FC7e#
/X<e6Re/-:IC,P4WE;gH)/&M+:6T6=GQcY]+aP[:ZdR/S\(II#e3Taf8>BSA1b_@
Y&D6W3M=4DfC<I4.O@BVT+A]]RdS<U[-;AZ&U?#AfG/M28fT?\5D[KG.b:<3a^RC
b.W_<5VTOggf.5OZYNY-^K\)Ng6dPASR1>#E8._fSB+A;;0M8c3E5c<;9cYG@)cK
_XS\_[7CPSO9/9#2.56(2?)faaDb::eKe33;^47@_9Vf)I2WR2\TRSF79e,U329>
&:J)NEIdT^O/YdK5QX1Z?&4/2GaKVTEG4IM9M3_-fWSd\DXKe/_-8CH;.9PL+=-b
)Z;S^b[U+:0Mb3.HG.[cG7EcL=C-7BQ@>BKI=;R^+UZVSUb?Ja9+6.)d\a,D-?_G
1KHPQ82Se)69[.SE?@7Q&50-2>L0R:8-M=D8/<M.<FCDMLH)2V\e<QAAK\:\RWgO
c=aYW)Pc+_Bb=@e1\,J\Yd&USL;a,ORCbI3=<E>B5HPFDO0:3K:WR&@CR;..e@:^
Rd_eTN<E,Q:OBXT0S>G:)5Dd&,EKB)]LF/4_&-.?/?/=:_3?(-)F?X3M,N56)H&f
N9W0eICN,5XCK54X@:GQJ7<8+@8W)0WYQ:RW=dPTYd<EOE?T/15X?V23]7-8Z#BW
g2=D33=Z#/[7f_d_E>=WNd&fKP(I70,fecPegTO]ZX(A\T#X@33C6.7I4AXb;DUR
#9MZLAZ)]EcP9AgCX;027IP2,VMU\cgZ.3B4VRSN,]\aa-fLc)c_8:=,GG5.Q/^@
KdC#D-JHfHHG2#]98.CgWBRA&^[S,Ib;L^<X>(^B_^?;CZ;Z#0ZK;0+MCCU0^)FO
#?e5>ZBI\ODQ-Mf+bK#V5>I(PMJJX@?W\1cP6PZ8U\[@(BO@:dW6[^\R]Z4fdY)S
LTF\eORIOQHL>YO_fI24@QQEdU(f]\1XKC;QQM8:Nb&?]WV&?H(@af@>O6B?2)0E
)R.HZ,NLSNVX3_3/U^aL\N+8)RJdOFOf;V.g<[,3>Yf?=gLOfS9f0XQX6<F\E#?2
3L-2@34?D#fC+&_H[ZGC2^1L6XbN.K55S^<BLVO-gUCRQBIW.,HW(N))QLYXLCNB
Y?YT/)FFX8+L);CbI5H^H9O:G=OBEIC31;U[??S3gaH[1PZf_O>6Fa7-;?XRX2,-
<cNZQW\EE9U/[:XeId(517W8J.RHHLR>E/8U#GD;6_=cST?6AXbP[.IW+1ICGIM3
Ka(#U[G6Z-08GW=0&<eE126F#=dd?b<PVDA>PbYcZb\S9Yc@-APBY?g;)-bI3/D-
9?<SS),M9Ta/TA.UgQ>5e#@L&):+3T\W?]_L\V(8f&KD:JQ^T)K-7\Y+-2A;eDNM
dgB@FaH87,([-@[:OV+>E@FH#+1J8NdZPC[@<]>7WI0-E47DcZBHBbJ8OU,(07(-
8=<eTFg7[fOHF0_#\PZd#Y]KO9)b;@^5:@I,2ZUX=MPD(&-A?0TT>R^9(,7^8cN&
T,40<B11;U?^I/K.[Oa6bcd>B&(;J0S-Q3cPP2T]]VFJ9f5;U,DQNFNgR58WfBU^
^TF;2O,GNN9c&BR])UPCfTJ#2<,OHRN0;8FN=?HGb^X->[L&.<b2=#[?UR>FI0f0
/]=5KWb-SJVa;X1W(Y&I?HTKD]K0,TJ:]055Q,#U6_;>II9S++(<Hd4P1=^(4H[I
/dGOV5<)a_f6.7H2e6Q4>4<LVXAB-=YP]+38WcXVXFM^bZ[CJ;ZYc,]VKKf2##BQ
dADF7GGLAKPNNdURf#2#RH#J]-J5&&:IaPddNDc\.X4#?/N[#<DBY8e/;PN5G9TB
:9[F[b])P>(a?aVN&3@38(DN/CIHIIGRA@4[/+TKe>XBTD(g:#4=F6HLY-V@A+2N
E.@Od#+EC0b3LaRUMO6:3V1NKb@@.)^R,??gB38=9X]bRN8-1eTL4]Xb:S;QeF[8
HGS^+ILC=ZI)@^&ZV,bFYUPCCKR7_@22O=ZZVNcZ9a09<5ZV^f5-Md8Td=ZX]8eW
&fL;2AC8/HW3=A#IRKdXP=LMC5aUfB6)#JIH[=a>2HVB0T1CCe_4/_9_TNGT1^)8
^<7Q,_/PXYd4]87STJ76fJQe0TE0I]LBL,=cUAb7\\6QcPL^)W)d./;78DE0/dL,
+?>L[QL]fO-fNGA#\AC:^E/&#<L;X]00G76](R28ac4B4dRKXNUA99aZ\D.-?ZYX
dCGgYQSLO_CPI^(GOWL4db2S/EFZVI4RXe5[M5XA?/9WX(50=+)9WJ/.I@=5^Af-
C-]1e_C1<f,6e6@_g:YeX0=V67>b>J:YZN8VJPX/b&E)#(.eB)T6Y.&TZF_)Q\fB
WO\1Mc],L)ZF&d6.9>acNN&-KaE(YgJ^):@6_fC]g3\@]gZS(UK=1+^X1XS^&XGK
CbW9BRa4L?^d8J,PM-ZI51U/J]gFOKVbF=?GbF2R,e<)+b0(_^UfET5.S;O6;X>Y
^6^\M]-DJ0T2d[2K[4HaTdNA6J#=F]I[C(M2QSBHea.;#5Q.RP9)[@EegLU5Ve?9
RFfU[FG6<+ZW42XWB8,+be&Y/RfdSd8(_&B6G3V],D3;Mb6WX)I4SI\Z2FOII6a(
#+7COD3?_.[Q70M-[L\E-BV##Ca)IRW)VYA?Q^)F]e1/RD9G[,E2DTd-4Jc=E?@K
<Z_JUEGd^V/Z:f@W]@WY53ScQT<RRcR\Q56R/\&Ea;FV7Ced6K=Tf0TQ4,-f57)@
?>e[(.-;V9##0eEgYeJLcNAY\bX\g@aIZ4M.3X@FZO7M6(4&.b/XeAGE,aM5MQ)7
g6:>(e7@1H0C>g,=/9\]D\]Kdae9Ka^Z+/VDZC&RB<:YFKMRE:D?,2)eKfF6B5,]
H0\HW<b</^,2^ZT+V_M+O])[>cP87;<[IF.427E.JTNNb>9T:S6gbA)QHS.HH6Y=
=d6&1IK42_KE50PZ]5:QEB;NP+cHLWRG+KA]F6-4U-):gJFOW0\/9:7F4(?L>7N_
4J2Y@aS1.:T,9b(-[#]=fGLA,[DM(b#<Q6D=KY/-A\V_X_\PJGAU+,9IA90A>#C_
N@Z(QGE,+9I-Y;YWVc7>=<CSHUEeIN/T]0G#8&YN-eVQ+ON;RcH,#01FVP_OG/])
@SHGOV<XF31bf^&:Tf;(bH/5C4F+DT_KT?R3>II]?TKO@H-DSE>G^1NL.VB0<IS9
?2#0fcdLYUGF4#>G0?4)JEC_C9+N@+5C09L\Y?&d&e3A@@GITO&=B8,F9bJ>H/7O
Ug3@HO@,7[IQ=3T<Ce<d-egb>Dg6UJ/#/g8+gVJO0YSXXJG&Y^VN61<5VCL]F1:M
<_,d\(1fM((RV(&V#Hb>E:YP7YS4GMHIDb[LS4>bV(g:9WCVd7Q->TV.=D^(ISW[
X,\G;^^;TUcV8CeHSd)d=63MB\,I;IY#)FeYKUEC1+@Xe+/:W--3fDc]HT<_^D@0
AB8T:YLC(Ma88#6gZ2RDaFKO5[b#c-_F3WCU3N@XMG@FL8L^]H5:a0IHG+HTSF2/
OY0IcI@FFKG<QG/fM.b7Y>T2TV[5@@ZK?OC^1LTSBO/aO[B,41&1W/34<@g5&ZI3
\-S)8T42.^c[:8WM&#LQcaOEZVI>\CWDH_;P9_JfLF.__SJ=/11d@1]Bg5_8ZZWd
eO>Ae1dD<+3-NU\M8TRgH2Qe4NSaf6(&RQNJQR8V#P&UW?Ie#_?3)2Ug>KEN^)IA
-+KPT_cT/RCD^+6?Nf[0Xe>ZME&07JVg56T=^7X1c6NOfFMAQ6e+@Z^Ueg+6=ILS
UN\)9KH0eOJ;>S=ZM1(e@,7e8JRUO]_94JS@#U?HI(QWI>9I/RS#.2dPR7-d:O26
4G?&FH7?0e3TMHKYY0dUJ#MAV(-C#:4ZbdFbG\S4Ia<WYA#(WL[QBT,0M;&;YM-R
3]9AE=^-d0O>3?H,CHg._X\L:8/>Ca-/L2JSC@OWR0[JcAB]cJ9BJ3-Td/fS;bF>
07b(JQ(.(K4^1YDO&WfTP]#U_eMU)Z6+e(5]3bV:55AQV6ZQcV1EX#\#eD=LT&g^
:(8.Uf8[UXW_Wa&]Y(=\g>S\DA#)1BNJMddPC5cFQ\R@]aa@596H/DNZDG0FLf6V
/9C6dRZAWIQ-0^MB]UgCWIUG8@PJOM;X-DO]K15JED@7\)2G=,D4851HCfaA1H/F
Z1(5)a-Q9A:bUa-&d4YD&>GY4=O1.8:GEZ#O&5KefGXcBHBRMg;@D6\&d0T):O<(
#Z?-9JS_><@LdTI@bbI0)@<ZdD^ZW3aH+g-[,1NF8K1I>5D:E;XX@(:[SNUDBZ<S
:9c44VFf^f0/Q(>7,PPWd_b.d[?b^&9A,J^PRPLaUE=5E6?4dfZ/]gF[YA[9R[UQ
V?Y/]6b>.Q.aJZ019S=<>2Z37<Y1F.FNLZJ7GW;aR#G(YAR:YOSRV0_TdNK#<+8;
3SMRQ<.B;O:_fRLN),4<M&K,7XR<X<DW-GYP<Mdd+;^\8F0eJD_2S@Q>L.48?H9J
;f?O#Z&HT>/8GcLO=[Fa6<>A_PKa464I8G+>@\7_RT#Se-cBY#>_FFbe5[)M2CB[
6,V-9ebHeO03g.]b0/-AFPFA^Oa19-L@6bAb7Y2L]&G4JF@ecUeED>eeREZF5#&d
L8c4T4J[c[.J<B8?dA]c)8-K]/VRN=&@a:.W<f>@S<LX)c.Y<dHPY]g]T#-cQ#B&
d_VF+TC]gHdL^E>)#RS<K.I7EcF(D0c2:g6-V=/f]8cP>((=V2eX(Qg>,NZ>2PCf
\+bOH?T)QW>QXHFNG0T#:E?]FJ8-P[=O4M+NGGJIFZY#/ID7Q)bB16.3SV382+I;
#E4J/.UBa+TRN@3TZ68HNU^^><)EBHc8bVR\[BSZ]\^dQ<P>EGB[gT2RLb7O&L9T
OK2V.#d:G3(?#9E7#M&B183_+DbCMeGeT1-HAEeb7PK/S@59CdG#U;XA[cMCd-N9
HWHg<[2LN^&6UAH_FJe6PRH+-VKWT]7^E.L@B##ba:&IU[SSYT21?-UBR3;e&Na>
_IKPe2=TdVcgDBUA<@FN(77BGMJd.aHRX?)a3>P2a#;cB-7#0=6@d>3d_5_Cd]8G
52b@G7V]2&gQ[cL0BO\OWUW<##d_cb]PZ06U:8cGQJP\O[^.>&1_#4O;2Y),GBgV
]U?/d4_#S^>+[:(HI^b\0-4ID/?ZgI;4H/433>H>-Mf(fXDdFGfZR+d57RD^7&^0
ZSX@<c[B7d8K/;SWJL6bR:W3_I(D5,-EXG&<(E<R7-W;31K/>C2e,]O2((\34L3X
g2XaA\A<+?W2HJ6G?&6;P;DI7M6,)3@TLRS5^[8aJGaMR\F8;EQ@4<J[H82NI@LU
5TH\N+@DQZTA-(e3T6LPY3]2D#R2PIfa:4+6X:L-J-7,?4S:SFPRV#K,>DaDeKCc
HR_<.F)?bA1[6f]P:89;,UM1Z5=,CR=4)@YGd,(@3TUe[#4K61D4H<DS-@QAV[31
-cTCeXNX#4Q,?@1A8GGW)TWI&85?dRT2W,RK);ed5=OG=4d43OWJ=9>f(aeH;??I
(-Q2RPOMbP3RW;)U8/@(AL(;O0\HV\6RPTd.b9/--G1=c2)DIJ@8b:&d#g,3fb<I
_?VGN_IWG#<-Yb9LD_C(&601\eN6],N5gcU(cVZWNQ,MPA<0g(]6bQ#Q@2E9:,V9
M@C8,-I3VJJW7A9R=^@6[=X&IMR9T\=DFV=-<C_:N6XT34HJF0,[)UGSM7GOJFYe
6DO,,?)EYe1U6fSXfYaRc@RELg0AX[ad.C_^0(_V?O(8:]ALPK/eHF,=P;QON6.S
P#Y#L8VeGX]\X13\T&&^7A7QO146R;+JOgb<WC179cRQPF-[_&.?)cQfaW>2^^.J
e=_&I_ANEZd=+B6M@7e<E1^e@T(\fD7abG74&G@2_gDU):/6\G1(faaSF6,]4RL0
]ZLD3]]M@3VJfdJLTf#/^<W+QV?CL7gg&&6KYIDWU[1Jac_&EL#?C65:#.Oa=G-_
&TT6_7^e5.^,<]@HK0,XQVdB6Z8BgU:TY-YcF]=:J/Y,7eP@+WbJ>.8K12NdRH?_
NaTC-W3&LPNQB#\8ac,FIWRB^#S/P]Y(GY@;]c?2K[K<\1d6<^QV,;7>\>aK?D;E
B&S=.24Z219e0.Z,,>,N@V;(R_=1\?]aI,1U(UYS<,I/aaSPbYgH\c:CD@4-B-L#
ZX;RA/a:,\N<LWMQ4\_LeYA_._<f;W<H:;]W;.bM<#MI:N)/41f0MD,S[@:]E7L1
Q:N78<fVT?;GDT\2G,VR(SKC(60(Sc\C:&?dJ93=[dXdKTc.1dVZ_4SXB@bXCC1@
/4c\][RB/&.,^O56Q6f+bg3aEE]Y<76J_)\[L:6(Z66K)^.\_CJP@G]ENBeHc:eB
-+N9TJKb.8Z7.W;.+00Wd3DE=F,KG]RNI_G2@RH;/f/+_NC,T&N3a9B:7]W6,@>.
X=bWbL\:S6W9\ZTe\A^;d)MATHP:a.B^+;dRdb(2g8=15&@_7T;cKc0aTbF^/,SN
cF6VFaG)RXa-VQ0=#eDKaA7\9fI38T)XaEaT^9J:MEc7.;Z04))WWQegO&R+EO_g
?_+16BZP+\\bfV;]@EFL&].151[J<C\4([+8X/COX_QK\QN>YO@PB(<TIZO&gU2g
8??9XY1g6E6WJW),Q2,Lg81[UfDd2WWRN(E9&.NRd=.3FI2A7PQ0dB][f28c4HaE
g]+P>g[TZ0ObEUAg6Fef84B.8:Jgb#^O&Db4/cW;8e^Xf@3BW)Z[@)7Y9>gNe,NI
d/XQ2);TgfCS_E:G<c=g8<@(:7&Y=P,,C8d?=8,C?[CRFb&Q_gT&#46^Z6?K]D<\
MP#(0H6UQY8=YcD1Od:^6ZZOS3ZX;PGIH,&N43P2,Q,G04HTW&Q&-d\^:.9IY<I]
A<(DV_WSH?.2?ZB)VELX3<ZI80GM9I\(?@FUEf175MMWA=2fXB.=HcC)=T;>H]Y;
/\Q7.Q4C^#eg08D(-9+&DCGIR(RW(LQM[c3+3FFHYDP[N-6Ge=g8+b98.RK4]\85
UWcg94DU0H<4Mc\R/#N9dQAC0\)OYP:#ZD@8H&1WWbK];9BDeI&@GJT(K@c[?QbM
PWbLbJFEH57W71:7UMaYEMS^Dg8NX8?Oa201K)AQGfa.f;0I&b+6I7g]M51egF?a
7Ja9A[KMa/6KE;X4O3VFZDLbQ&cLEeU]F)YP:AIf@5M=:9]POLNS;NBWLO2\LcCN
A^R@U9e6^,#gINGB>VLKST\>PW^\Q&O#eY:[fT7/#ASfAMFGHaFA2TZ\K^Hba/Va
,GP22_(>;@ScFOZ40CZKB>:.IYF^N)M)K905&B36_)]PD=J@P>d7g8)Y2DS?)CaV
7c=?7=AU_g<Rd5;Y&(:>.9g&8]Vb.7\U-2^UI9XaJOd-#=^KA._V]SF^6MTHS(BH
ZU5J)g6A(Z)BCW]/WV&e\bC+_W-0PO3)c6VS6bELWf4A;1R\M-GEaf<dUZ>48UY\
c78#Uc(e1.)UGe&c=@-./5[,BX>cCOWJCZ&OY_CcV=d_NJgHbW7H(^Gfd8TG-E3Y
^Z11X93,S9Y[P[TWQ]Y,#CW0GRP=I;X\f]bE()4f4<15QgEgI5dEfD@</=]:e-)R
K7>52<EF.#K?RP48@4bBRBU.BZ47]2:6]QPU]Q<bE1?62_W^+B/_><CGU=MD9F_8
1XT:g>TI:[d-Q;U6ga5=GUaD@;/OeJ&-<<afWD.EWQ<TEA(Ye;b+.)>dI>E7654>
>+&U:Y),0bRPQFIM9U_<3N5gMVa;^[f]E@8abJ@V2d84IF?GaD3c4:6I+W(2U6ed
,;Lg+S#]aLK#NO_CbEQd6&#2T26_9FWQHQT7=IW[Ja?LSYg/_-L]B)4fQRY-ZfV9
]5A.>^7gXQCaPU>-H-56eH8WP<De=F&@Eb]E?>Yb;+40)1<Q2O-5I1.B-(^9_@:@
KfB\7K=-+/X-CK:_\9CEA4TaCf\Z4CFAa3/WBgg^GaW3RC[:BI5ROcQ?[<-F-RB.
O<1-W4ZdM+RSO\:C/DK[fK/?VMff7[(&f0T&0LJ:+.b>.Ba0SM_JH8>f5VEOd7O-
;QY)L6R#Hd5#^N=@La[SUcg8bd4@,eFY7L9Y[EST0QV/J;J5@Y>?O+M9\4^+=g_;
^-=QgD.O:gO:R)1]GY^,a)PK^[BQ4)3cOXHG[5:;-]Cg^<;.B@\NTDBg6[N2<\@,
DRPWRDQ?2Fe;eKL,edA&#BP11UDg@S)Scbf&L3_GW+a4_:R4K50.d,(]O@.8XQDN
E@?YEQd&X&WP/d8(#:J#,AZK_dL)IR=(0Uf+:/S4U[Y6R-NfK(BCV+)4:UefB_JG
Pf2@UI[S1/a#D_ecfbH&UPZge+6<,[M(O9G=I68HI0+ddf2OV0S[ZTT@+X+TgTEX
-9<>IPbJ[.5)gFb&YfMMND6c<;YZg.0VA)[a^]YNHeUT&?B(_,b0D;dOdDH2T9X5
LQg6b?O4cC3>+Y8R[O@2F^<U5Q5O@5CGCQ@32KY__9^27b?,/MFR:;bHY_;W-M[Q
IO(a5,<?&b27UUJ2:YGHe[H.[TO&&C0aJ/9f/J:2\W1F488E83>VJCPLKS+FPGd:
XD(G6b^@Kb/5[4QGH8CM=/YKB-[,+?6E[EVf0?\JeaJ@FSfaX@YR8)/W/Z01)E.2
:)ZU-2G)U9L2BZ]f5T0#H.\-);98PZ5,J=G@DIVWN,J=6[/->WL?c=_=CDL0e^0A
-&;b.cW86NJTdcfKNL1/Ud.I(CKJE@:T=YaXYgdSYf?=MNG9TP]f(d/&GS,TXGKC
PHBA7S-;B4BB[@F+Bd=>F=e6[,Z7)XO0gdU+EFGN=@c);Q)0@L-A1]KQ?4A:-gD;
37V-KW<Z_.fQH\=6.B(>8;c_=9=1cGa&[=aZ2Rda1?MS>D<O&?)Y4ffK?a(NGB8Z
C@:@@;]50>gKB/GHE/\eKaB3QD;d1(KT^5:JF-;,D.NJKD#.O<6Mf-^^U9DVF;T/
fP==.Q^@?+#2gY;C^85),A_KabdgLB](/P5(.ISLgLY7+QV?5fF:E2d#,DU;GY0Y
.dR2ZTHgb-4_Q-Y#WF^^3KX.WKCYG4Rg8U/cf\@PMf&T.656ZTB]C@GC?Zc/db\a
\Ne8;@5Y(]aAf@gNK_--fHGV,U)US2\:5D/YTJ^SB/1>G#d?X-[/g8A,7aG_:>M8
]G5\?WTPT./gBLSf\;YeC+fL4^GbMFF6bQ4V-dVB6VL./S3DO2J_DFfd-H_P3WQL
eL]>48<N(gCRdT@Ud1;:=@+2MEce\1d87(UASQ?Wc)&RO2<dN#2W(9CL9P:HQU6A
fB<JNfG#BNND7c.[&Y;<:@9X-c-,B)D>ZDdZ)HOfTLCeP\RKB5+1b:KXU9UGVAWA
Q[a^<XV_eUK\\Z6IJWL3Q++TE50QB5A]2J+/2-B^\:418R<W\8U6WZI_Af__(fcM
@dgEg];eUV6TZ+E<FF+)^P@d5Z+SINIeITY0Qb)^D)-_L^,1TDY&Wa_J-(aEW04G
_ZIfdNb8BOcZ?<KNf(A\8K&I,bd86Q#]2b:5P<TNd/?V7PH2W_19Z6;;A9NNB,25
.3cKQS+1D=^=1f(-E&NU4c&/^C70P#Z2IN&\.RB4:ST9#53K2ab2NFD0a)=ARWP.
T8Y;<c(<^3B)L:eUcf4AcI=aCDJTcY>Za=H0:03J:\_7>aKZ\c810.AO/N_-8<Z=
:/Sc@B,B::(HFfAX8>OP7J1ZFIF4ggVBVI=J(X_b#b@>;Z&DZN^]PV^M:\LE]&-A
\eFPbD:;O1]XV)L\#+e@g351^#&eAdG>XZK2]cO@^@If8..)#e;M5UXVaX58CF]F
eHT/9e-OJaHK6a)6gH&?@\+LPW?)EI^89cX2\8,R/>.Q--V@&K8;HO#3)6Zd<>H2
ZI8KD\X5U[=96-&X,\6CY6HIOQ)G0+2NY7<9;V,4S)09d5UM6^D#JT6@f\R&=AYT
&5IgL8^YRBMG/T)HM+;;eW3E[M?;9#-?NZ9CL<O/T+]9MX]f[,-J4\GZ8C\\TdSA
J]3DAAdOWf[>eS#)&95PW.M4bKNK;;;\Y\X[@><6JcO2CdFc6XL9Ndd)J3P.2SV[
ZIYKaTc([-/IWbQTRZ0CB,NP6H1AA4A+C,Y,#?V):P4@S(9W\dN8eFYQ>>TB51AD
RYLG2,-[=^bDI(Fg[/\_>c>#0c7<KTAaE<>]:OH#LH?edW\IGQLWV5DQ^Ka2G^V(
(1B,N09A1Y?H0\#4R\?cfYJeC(NeHUR2<^OPAX0B5M4EcCT)C=^JS\G07\1P:E.7
bZAP-BdX2&QFMD\WP;&a9FM6QAg6[=>O3c-[gANg2>+\8FAC5K_\]0\QG0W_574N
H(V&Rb^61LFMa(]Re&7:,DB&ag\ND9HZbg+HYf#YUY]GZ;X3KA<\>6__^-]\VLO)
QNWgEF.OJ-BE?:SfB3HDL=1&>9)B4X<<8,g_U<V:S#-?R+TIO[:1^(4-8S-89HQ=
TgHNd<3NCBM,Vg=6V^7Ud]6YDg-f_M]LT/>+gC;T#UB[6IO<L7G+.QU:ePMN-MM#
.H1HC<\B+B#.8ebZ=G<DeVRG+((&26g>LS_BT\R/8#Z-?&S.@(?bfG4/dcHPM7HD
B0J@&^-T<UMg:0VTdYOQQ(Z+ca+[@)b-US-DJ&Z>Q-+1CCBZWcHG=aW3_EFFb\9=
^/M[S2&bcZ3QUPVc7FC:@N/^K]?7:XbV4JEX/<QNf@C[\;cBN0;=.]+bg/2\5K./
M9A2X<N^,H:=:BU#;G0S^@^DV<ZWUW:3=WGLB\bAFZI\H,@::&OY67J/KEIGLHC(
15GBdS(+=,>=B8#g_+K7B;<V_O97>,14-0cZ\?fZY\,U0SHPE(+N5/<)T59>+C_g
0;#c6:^7Od(8F_-e(?J>Y<UEVM\,^A0#=Y7&e9KB5:=GM=X/dCM]6TR0]P74#f5Z
;V(4H+3(/S5TGeZ\<#3,Q&+W8FD8/AEOE0PFM_G=OPYF].Pc:GW+.\[XD^O]M#]\
VT8AP(0]PLZ,Z0R\c;00<>F:E^:7IS[B#=ZZc:17[#Ee[Kb(Z\[dafM;9g/b@,@(
1X7Ha^]92E6FCXG6TEJWHOS8c=GA?OQ7Z@F2GcT\,cB_RL=(PKM9TS=6IR=X@-\e
e_b(YCP#b]#H/\I79Oc+E:a1TI48VObJ9-TJ<TN12.T^.O2b)ea_PfGNVPJI>fLg
&8<H1DK>,:@aJS_E;7RQU;^X/&<0YH@F4,]\7Tf[aY^;SN94M4[gK,QLE3MYNW#,
GNA(d\AO7,\fbcO#9SGKO1<e9[Y[OZ\6ba>QP0>(0;CS_KGPMVC8GKf[D84a8IM7
F[V7Fe0RcCIYd>8155/E_IW41&?/LIS;F5;c[LW<&@.ENCO)L7b]&ccNSB0c^C5&
RTUMX2?\?_A1f/eK<FI\Y#TR?aB/+4H/(bS86Q(<JK#c\Z[^RV][/<<<]W7AI1:?
X>eS[[e;=ME;?IG>H7SA?=6-LZIaFLbW/A=Ea\F;CA+MO@#^QINa-If^=e#9G5?^
01Qb]cE@WObfVA6T(aUa/4@8CP^:V9?FDB:29bf5\?I9A<1\IeGBaS-[5N\eS[-@
J,KV^6,Ida@d4BCN_BfOCcP@L6QAR9?Da&(Rd5.AD.4/bWN]CRYO.^<(J((I9U8?
Vb#d((ISI<^^UK.(8OeMK93SS^a\^J,MAgBI_=#&b+^6Cf7Z+OGSGQFX+6@UB69R
]CUJVGKa[RgdUdDON9#7(ef1,.4E3D7_>\RNL2DI^V^_2O)<_)OF&Q/76)aJ-XA2
3Idd2_KZ1FNX&EDR9TB-L7-818W>,&f16YK(]@@g@^feeS)13+4+]KOYZ<B167OD
LW.U4d]D[L4KCNZ7FXN+OI9/fZ/PJK]b74;QWCV>\8H,Kg=\NQ,T8:.^SAW@2\;&
5Q3:Z/U=AT[QUKMKOg95SFJ4(0.#L/Cf;(U,3g@39W-?3f.906V7+N#,fRO-M59a
S64,WZWV,WFS@R@2(;5RX.HDO5QG_G?V+EWM]H&6J1QgX\UG+[M6gD,&3/]T-YN/
GM1CAB;>aY^eH)WEF/LfP4KDcUdWBN36c7=(bGT^2>T,,P_8Rd:He8@cXA3N&V_N
7LBEJLCcBdBOYHCWbB51FWWSAe,?d>(2^UTRE5SOWYK6LSg;,^c>-[&L7Z0BVZAM
C,)W95/^bMc,gIeD2HN)Q4JL^_R.E5b_<U>)[(8L,Wa5VaNU^76_GEXRO83F=e:T
4DOSGOZ1/5I]3LDK9]QfeQ7CH.)+P-P0.K:S)@IT^PSQVJ3BLFQ96@O5Cg/]UC>>
S(_)&P>0N-#185<1\-R1X>B47UHOc].:Z6UUI679]e</1e&8J7L5VSd)H62FKU7G
L6KQPb/AC6<&gA?L9PBZ8#;J19aJ,6-I@-NZAB7.)cc_NaT>ZBeJAVd#/:@8]dgV
1[B4:<C_9_NIb3D>c3D<Z7&RUTD0VW\]5?UBT^(3,/>1]M5?fU-,[[;OY_ZN-?@f
(\M+JQc(SfI\@4K<UJL9Bg[D.\gBLF:fFW_R7^d;R<(EH1,;O6a]B<&,e]_0eRKD
/86F,A\PTA<d\4f)@a\:0+A444/J+#1WZLd;VJ47^A7K]<J0)&DYL#<0XIF]efF^
>eYd^S5_8.FH6M41ab5)FO<W_e@N]OM3dE.Y3e]TKJ1<ST0K^?)?VQ_f69OFFDR,
,9.V,g0Q3S7TRO9WXC\P:,_^IOZcb5Cf/fCN(C91_Z.aW5#F<+/+G6I2_a8LE?eS
AH<a>>[\\7F5#<.AA23eMN46ZLeOeSZ:J/=/3Bf01^d-PPcG-P07#K)EL>_@M:TG
RZFPaW5SBXO?HH[>)/LVSf5=:0J.TH2.f/VI-G0dHF;_373TYY:&e[gPG&Y-?J/[
M;8cD</LCREA-<9.AFL\Y@.R:,D)3<L-IDaW9:1eV[O>919a0F#ZMK^=#ca?)]Hc
P]G4WJ+9(/4A+gCe._?;TTd2S7d2a2BL>K1(38^g6HYDD/b2aE&;L&YSgN^^=-1K
LIW^A@/6c)L^ET;]=)g]D^(UG+C0.8J&CEd1M4a,aHJBKa?e[.ZBd,_1McO8fCg3
N_7VdL@VZS[SN]fKa,?RP[\fA.Y:V6WUf?aF]S7?V1]RdG^?^-GeYWa5H@//_Vb\
3N[3ZAZG6(6E/;;94WX5-&FP0RWB8,JB>^EBJ:b<Qe.K;<96L-1=c2F+ZaQe.:U[
QDRMa]Rb:8OWYY68e3AGF0cZ52@]KR=<;OCAQ@KX4EL1/_C?7<JOB(FAg8L\M8,3
VV\4<.-f@GPUCD-&fS>DW0f)_&H]D-bU]2IDeQJR_R&7^S8GGJRIb1Q@T5R]cT/Y
EO6X48)@Gf=bd-(?UEaG9BZ=7;EC]6M(ZIY@bC[VVFNNU]O6b5+IbEJ\N=dKX&9Q
dFW0Ra\[94VU3,USK[R)8GHG3Z6_KT&.8Bf7Q/^SGD[,MA?^7T)<E8C6SCTNDE3V
8Zf2+=16T26D1=C65CUWG=CZVQ<?ae#?^\0+=RBUPOgGJaW_H)S_5>Y2>60LUdHU
EDK,f+[\16:;?:Y4USaF@&K8OZ6B.P;H6=bLGK/[<6(^;L.O^?&:@NM4\T,Vf6I[
7+](JX98\FW=GdBAXG55e^Pc.82NB88b[0EXRC)(E-UG[+>(#8>Q?7UI:2VG?PL3
5459?T:SMO?#>STF2DP6#9X)7BP@&K^C/MK:TWVV:O^Y^_7Ub]A,]f/:DFeZ.9KP
0A[^>Ig-ZRX><Ib-:LPgQP,Sg\Ug:0H3\Ua49,]?;H7M(dcF/S6((D_5R,_ScS-A
Y??cXbG_157HM-=;bX4E;F_f3W[+(&d\[X7]++FF[P/55JYT23CQ01]E\YQ-3#]/
S#7ee&2/\#Q__Q.&=<#(AH..]Nd),(#NPW+GE-97Mfg)E?4#g7^);E1\_O=[4L^^
Q&NXU);&2M;\EP:)3\Ce_T9Ia+=.[Q>4(.d-aXdOLT9,VSVK>>K+Y86A2E;JL-Sf
0-XXTVR6/T7B\-^BZ&#9H(2Lf#MRg()GMd/fc-1]GU1eaEOY5c@WX8<?=MMX)JB;
XYISa+6^X>U+B8\AFeUHBQWfFAWZ9<]g\&,A@USa@HI<I=CM&JL=cM>]cB4=F0P>
V1Q&Lf8)?[NTKG+,JTU]d^HaH34N>\,7;G(<@.1g_?IJeA5T84(N,RO/T?9Pfeag
VBVGeM2Z_[gFB&//f<OM9S^@G=1Mc;&[@aNH0U.3NRN9B27QA3cXJW.a(E02fd_a
@K;4cC9M76CPKBKW@&O32c2DS_36I:ID9@0;LV<3O<?A]>XB>J0BO30LC3+CK)I0
Yg=;(MZXQ>>#1ecR3@,g40<<>cB;IeD,+7O=)N4,VE+,/2U^#W(S#&QX8?eLb=,@
IC^-<TQ\90)<g-Uf^,b<2YXN=^CW55L9\3?U4PQSM2E&YV#N:W:FJO&L]P^I6Y1Y
<SeWP0E<MN2&TWAR?+3a6[M0WZ^KBU>9R:&IgZUG>G?OSJ=5TSf,Y3B@-\M+&cM8
US=d;B=FX@H&1ODINV9YXIA:CO_P9e?3c6bVb#=YD/PHL]#&1Pc#,dV,W(.,FI85
DVKLGCCX#+[M7bT812FZZA>8VDEb^(773:8YT#J;[E\JIPXbD\,@<AQY2f(XXMJJ
#8.e6/;3(H,Q>TY2]P33XJC1HWeCd7Eg]e9P@Y5?d6UL?0W+@[3C#,gd(6gfGKO,
[/ZN82>V;73<Nd7J,DEdLeRPgIO^f=B>HH5T,BcZDE/_4?^Gb>K#M=g<.5gYW[.Q
I/d(D4cE1Z:b4:)LTPXA@1HM4#NF#+aWYF4Xf?OCE;^0dYRa:(ABOIfMTDPM)#>M
B>.-RPF]@7QF4XU5Vb_eU_U;V.f0_EOUHe3HfZ[?c0KB3.Ng:IJV_AQJ:8UE@FaY
g-IMZ[A/>V2GB8&?^fICP8\c](DG:]bV1JI(Q2QT,X#,CH)gOM:f8S#g]>QcR\5N
;8Q9c.Q(4)<[c)#_8I#K]<<#V,d>SX<\gZY\[fZXK-aY\+HBX[B?g?aD@P@a\Q)Z
12Cf^SH(4H@48GI([-/C#+^2-:5e@&Z0;>bfYPFABDLMWfTABFB(/4Pe>FR3VUe6
dD)GZFdFaaBE#FW3f.ZPXY7-PGWeg&/__VX]F.+4HgC<?2(.WCdad][d]-IY.==,
TO)0H1CDTKBKZ?ag9VD6AX=[gCS70IEFJg25g3dWJ<&6A?<A:aK3W-\cB5E4Z7YG
C??1\g(&T9)J/KGQefQ+ZF4.==DQ=Z\2I1^L,EKE0U;D_g:[R>DQ(F#W&;R_T/gW
AC?H0S,;S?J=8\),a7Tg\+9BgeXN^S_?5I(\I85DT/0dQQ_BdG0Z,+8N4N/a#Zd2
IRV=,95L&JOTFCM9d=I)YDE)RgZ@+gbK3;7RF9H.L[=.CS.>LC_J2^+1,A@_AJT6
EXLE6RHE]a[0RS_PZ4#M(5eF1J@Wc_/51760deK_G-QQg\3V9K\WcRf0;/K3NTg/
#90GdHYE;ZOP-W5d&.78&/XR,M632fVA_IEgI<>&])_IAM?f_Aa)?gIPV?QH4M>T
1eB16)9Uc_:g2?:6JATd@7243HZBH_aRdaM7)>6gDF6S+.(Sd.G/e4P-:.?BZX;Q
5WO-Z]&I?;HN&=:[.+HOFZa#E1PedS._1O<ZQ=A4YI5V^V4LZ\eFW,\V,-(R)dY7
&XC?@5WeYMg61:29FI;SM#4E+&:X20PFJL:g(QWfT:91B:L8>;=.=9,7\P?.6MWa
5?I#[12#IR.&IfT)S?.Tge\BA1S+Ra&78Q9(9/:>R-M4UJO=f?6-4)3Y(I\aZEgN
8WXAc_PN^6\C1gFWHIC?;eFAN4\f\X-VSS85VcEU(:>-Z-HZZVDWdagSS=9D95Qf
3B3\;1)P:QZ]&;2+F6R8([J;]Fb[R-Q\=NA0_>&\Lb,S)0OUK79N[=HS[ZB\PP8H
g.OeCV622-FccFL2a0=cWZPQ&?IC3e(IB,HHYEeVa_VT3<gEKK-SW8(6[R5125L3
NPK7_<[M<TJCTb\e4^LgFSBb#2:\)L?<)S2\6Vf_cXR/=#JD/,389G0UNOYQFbPY
,fPBKa5UAG&N_0a6eTW+KBKT]I2B.[WFC<OYe3RN,E]2a]F-WW5O392Z&E8C#7d>
I]N,Y##>1N2TODIBCB8W=&U1]PNC=f/-g1TT3T/AJ&C^RU3S020&N=I@2dVPN2,3
X=5N2b?fA8)R?OEL^N>HB?4V-.P@_d2M8R4T:B451>?9:UW0MdDGJGbN=HU].fDa
H=Y3a(YgdVc9gdEA[>Hc57(>IV&ZN:RIAEFW\<=@5VHAV:_WDO\b]8g0H&>]T7Te
HOQJbN<2GISWULX1>J9<?1)3X5BJPRN(UKVLU;I)N_=6#NH=7QH3g>ZR2F2^D3S5
8GODV<YQ(d>^=W_S>)L5#25<##YIP(2J^@2._?Xg=/2T]T&,W/DX0GZ]<B44BF=7
=gH>c(:I>].<<PGS43@O/I#A&eC;b#HdVcS5-QCbG>aKd2,RJSM5,+RERZJda[2B
6c:eL_PMBEgZ69U-;a#9#D+V1=fA@d<WYTHJ8WUA(+a+#Ec14PN<1>;J7Dg1]=#1
K_.LeZ1Yb\G7]g1g9Ne3QNW&>L9bI/=&IT.MS]ERC/+^>NWRO3KUGX;.G)NU,+2>
1eB\LZNQZP+,Y(KHUD@EYf-bJ#cN-B.=?[,&Gbg46=D#2V5bNgI6NG2/MFRZ-.N+
\F5LA4d42T@?KZ4B[0IBTRG-93:D.]:e:\4,3\0F:S9T^P&\Q5SH(;;P^?9aGN;S
226(baW-&A3g3>I7<N8Z=,4cC+(VZC&]eURLNcdgLU8)(>eI&1B[gcF#Ke[)#0&3
YD#OG>71+LCV5X;@>7#HJOTK]8=8BZDMFO54Q,]F>,;6C@LA4_UAgWUG62c&,BK_
OaFDbAFg-f#B]]<PYEIbTX:\;M(1U-#65::[OXN99>23VU&Gc(0-TNZJ>F-:;X:T
3=&KeRKX;BA1XSBJ4Lce7]DdEUOEeU?7HB#/_J+&<<cK,K=W&8J7YFLPQBCJ3(^9
7C_M_/V9@QDb^NOHDH;25]C0DIW2+QF>5U7]RaOd-;M&fWE)LAd7dXGM=L(GR3g@
5=]G;#N+[,XK/<+/HHIdKDU@?R1PG-3A==bC(^4Z<\6f=^M9S9.:HO:]N0e-8MD^
/L=U#=+d)bTZM2ERMG7INTH51=KR<J?-[/A9OLW9&g3@AfG>Cc]HR_XX2FEF+0a6
G7-gf>G_],dLG7:-M:K^L1O2;6^H7U<DGD4UB,gR-;S8F(_EMX;VE9ge_IR+\O0X
F/MFZ9AA<+[-HVJaR0E4g5VDZ2SGZAPZEAU01Y0[aPK<_<>,aR@3L6>#-0^5a=X.
cHIddWC@HX92245.>c0^M&HHDae[2RSS4OA:_]B7?;Tb)402\]74AW_a,+JJACJ@
CB9IE@4-]a.C\O]O=@/V-XOXI</30SgV2#aYgdKAH6WKeYG9HV]]F+L2S\<H@OKG
V.+67=?ED-R+a\\OUVB&/X,PgTF\OTPLGV&e1T][dWZ;P4OHQXdK_9f[G/#\bae8
FUBC:A.6KCd4)M8\0f8>Ng6M=R/R4\+aIZBOOPQ)Y^8Q(Ub5TL#D4/aYZMeU:b[;
I:0R&UNcVO.7TR.IQGNH,@1&;:FOG(/EN5RV@X&@L9fE/D@G2-/UL[?edXIaQ8A[
_JPCf@P1-f[.5YX7VIg&WMDa_LMEP615:#ECfN):bS.^)L1V+eDY<53?5d4]f_)\
Z=G+C&RXe6_Q?52acE_<1DdPIF<(J<L,JM.=#<CB^Uc77UJE9206Y:/ICMSJP1V;
)Nb7X8^#J9]:+Y/YC](GNAAFf>Jc3Rc5^b-H[P9JPfc7(3Bc0T?ScSXC?6<SM:aA
Ia+[ZSR9T0P5-7/gG#Y,T._2I:6V]-+eS;F@WJCTT:Z=/=fOE;Y(;IO;F/4M2-:&
:+H&Ye_Q.K#\:(<;PZL_bZ7;Ug].&32bV)^cQHT.BX0(>W=@X^dO4gBR1U:)fR_K
098b?MR@53K<aE93O3U11]0UF/;IU27g[E3(>d=3.06C(T<eHF0IS<E6X786e11Z
+J^<M4CSbR9_)3.SJ3.+fa;bU1#XF=U9K;8:Z]0,]YW2#H7/RQ,T<gVM6PP6;61M
6EY2Y_FD>EOQ-=2)6P#/5NM\Z3.K+\7D&Pb_>KN=T=YLJc>R?g/MU(3GBccVIad;
HJE?696JW;@)a=V]b2XX9CR<Q(]NP:b9],?83<2>d&2&G;a<6_ASL:g)gP8.N3)M
ZG571W>F(GERYbW0.3.JX]L/O\I,_<fF&>3g:,Xg]0>DZc]88I74/U3Y:/27CR[K
P(aWY\^5?EgHWBdZ_fW<\0<;W@;OJQT9L6VV+8)3];6VTHG.EY:W;K)Q<f1MSDeB
:UP+K@:G3?7:gF\c=_[gf+,A^H5-_[VdJP+a+[;?7X)AX))P<X/cTJPe=LJ7VJ2?
gTSY30^/9:5K;a?T3U^EIfa+W&#b+67\6/[0Zb69LB4XW\ST:CFC.I5XNc;:7Y6\
_4@c(G0FF^_P;<LaH(?6MT95MLKMQFW0+d?-LM:B85\CFbEE#:.Z3]^P^QZ&K].g
fcSEUI#aYZIT5=;6S1]P.b(<[K\C[NbP7CP09R(9Y;_F,:NaNRH4HLSR/<-/f8>X
NR=<d8X#3eUA.JA4D[M:9N0E-^)ZLT)IF-RK1D3LfWNZ&MDS;[O;)ffSFON8&;_2
aYHA.T&Pdg858.,U\b2^\dgPKQI.b2R(b0fDK>N<@;e8A(YNRGJJTb:>Sc>J5B)M
G-JYZ.)\@F@).Q4DYV#_#fcBB/,SOQ<XEU.XO1]N(WJQg[_TgAWfD2g>9BML4JK2
:]+87BW&0,f&d+4J+Q(bdcI8Oa:),9f&HG<Pc1,DIU<_ZELF;-Q).O?f6@FF>1BE
<0)b1g)KbG67_C<I&<)IcQ2@#8>W=)aP-?dM0<+T0?GL(bAE_BD2N)7TUa?(&c46
3Ga#NZ)c/P4O;)C&#TeH;[e(@H052G^:.8QX4T#,)@20b\L:^GcFdODAecM,/_EK
-L=/T;,&>f_D\3Q)+.RW?RG@H0QgO+RQ;QLZCY83:4aK6_CN&G3fUB&^Y\W8,:?#
g&DDgZSJ(#)f:[-^ATcbT#cP8_EbRGAf4SZT>HQ4/fY:aB6fN@5;Bag4[dAagL7;
:0725b+0NRbNXfN7>)SQI&)L[A[dW./-?#=YK1UQ:EOQ2UCJe<]g/<J1K(&&_c,Q
QQgb@BBKHBAa4D8:JLW>#G?=f8-+[QP+]-6F=d\bY/P<I1K5#.&(&EM13MdTG#8-
>JCMH#-:H>SVWZ&8XE6,,HeM7C)UgJ-J<7&[\eEW3ET&;)Y2XXc4X;.c])MSVf+a
WUffQ3]AP=g;7M7:+dSgKfOf=2:U\(\]gY9b)8[U/K(E8Ge>5]X<PL?a#GZAf^UE
L0JG>?Td14,D][1EAV1BUM3[cSZ]9ZgTc-#+3MG,/QO&T[)38Ed95SL;c0LI^0GW
Wd^g><MK-YB)7&c#C8AVXb0CW5-RP:X[64UY<@-^g&G09?=)TH+#\WJ#;98F5/ZC
@[W8-5+bI#-1?D+Z?QNOUASHC:g2cCHVLU9b&B-.HK3ZN5]NQ745)WPQ8:^P,:/K
DV/)^+(9685gVNeKRMbA2aYCdP.+5BSTaL^;B+9_YfO2-G+<#g5G=XeL11Cg]aQ@
ZKRA13TZ_/W#6#<,_Y=Mg=>Be-IDb.3Ad4F4:MJa9@E,.\-[W^H&7?c0BX)UbPEN
5==2+7JDL]^J:+M\I/c=L4]O1<=b[Bg+Z\0VSKBJP=M3E&Pd2FBBL^O?]<>Qb]:K
Yd>2Y/\>ADVB3HJe1_SO&/)\,0P-2dP]Ef22X?#U4ffTOe/QKM_/:Z&[?H@HX#OR
9P]#O7>(&-2/N\R[/TE?Eb1NM,M,<MLFM6#U\Mgc01ZK/6Y:0Y6[c;R>]=R4/):Z
<7GH2D8A_2VdCL[Q9#.PNRK;b0BM=&^YNL43ff5M?^;4BeB6(:gNd7WYHeIUYMH_
\+>SOP>F=G6F^9KPf6#(f;S4f1_Zc)-]#DbEM@L;3bX&-aSaQN+@)]>CF5@+a2d.
Hb+dHMaNP@>W/g&JF1_^GPdIJB]U+SNA-S6gZR97-?g@=YI6R][3T:._[3+2G#+I
[M,D#64ffH-PPD1:EX?4K5M\DV3_NKRV_0/UN>D4Da4(F0Q+01Y+BCP9-#5F+FR3
-9Ea[.TGC8^6?eHO;9DdY+Wd1@__/<D+&LIAfFf+=ZJEfddG+\R(:K1.a:G.0e]B
L4-5B_eO[DfAT0W^=8R&?GTGTd)-9X#Ne[CFS.40Z9FU#]X4,T-2a_#[)QWHN7VY
(]A+P7J#=I-La;O8.S=F,7.e6+-V30S#R0UL^>5/H].L4]e^cN0@a4HN)4A)4=WK
>2S-ZZ<?\RJ@L\\XNIV?VeAP1<E)-H755)@OIBb@(BFAgfM7=0-DJ(UD=+&<;/W7
9(TcDZ5HVJ\SS/3:7)YW?fT0+6HQXPDgT3CUE;8CO6ILb)f5T9F78JP)9/U6HL-=
/J+W3A-PXdZ[Ve?70^A(EFP.I3UT/?>)=W&(.Qe#[UegZMLd9C/b;RNPKRfZ:30D
I]C)=5+;34XTF1=YHU\Kg&cZFWD.GWZ/+O=DJ]K>;8JT-#d_[9JFT)g@1I\#W0c:
a=1:@A0NWJ>MB++?NcffOYF1^6V+2T3UPZ6+@(^/6\aF+PF/>Z5bNfP5W[N]a+=&
+-<Ced5WLO>1?7Mg,K6O[R:YQ_PEI[(>&V/e[=_=^6B[8IY5F_0Q2]&4cbQG3c9\
Ke0ZNDD?_>?6,_C:=)]HMS4eZeO<NHYO/Lf-NJ(CT;\,cZZ4>DPE:P_J?7>Z7]2b
Pe)aRIUD,GXB0Kb<Y/B<;cB^VH(0\cB5Q?Y=_HW+YT-U3#REDINGLUASFUN-2+F.
?X.4dbW(@;DK>;#Nc2/-<:U\=MAB6FF]P9:SDJ8cR;e+40Z8VL:I:\[VfC;PYBLc
MD.J4g8Q?-LbZY]TRU\_&YNegdQ:d@/f31a\G&T-]M]WXI-]REV@1aZFS7([MX]Q
<b5O+.O??6VAP&:_XJ&6-C)^&23=/LBZO9COCRJ76Z&=WAZRF^,PGN<08M01<)g7
=[B8R>aJ,.J6+e5IZ6#?#_3GL[YYU(IUHYdQAM)aLM\/ADQ[THSAIL]S^/V&5=)P
FSJAZ6[?@FT?5a:d]>MD&\?Y>R7-#6DJ0OJXFQNKda8\JIB^_40=00Lb69\<a7:M
PHIO(<CH@fP6E?MScKXCN0O:KAJZc(,e>_[Q_.E0\D++LYbaKBcc-/)cAF46517b
SB0_f92OGcZ9aV<g9:[:<Lb<PUEXIdU.K-?ZV>G+f\1]#;21fW9d0ZGf:^WUH,=V
.Aef_V62eQQXIXH3CI[(g<G4aJDDTLC#UTUJ5g+J+_D,e;^5LIYP;U_=Q:NPC2;4
^K@bb=fXgZ5Q<Z@=b,]42HaTF1Nfb6=AE,XU:5AYKGB//OM#XMW>-O1aYBJK,1W0
[>d9MZN(5E&4e#O6GTg&@<WB1H:X6X1P>/15U0Ld&9-D_TPK4_+FCJe3FCE3fPWY
#(deLEOaZOd-&2eC\2[F6YI,MQP^4gLG@D;@-Bb1X2_7>R&:b.[#b990WdP52OE\
aYb@db265c<9Ad?,5L(9^Z-:BLJI^P4XeV-?<dcS0<Lg7XPf(VQbdU=JF,\X?B;N
@aAVL,)-:XYD=eF/a1f]HeFDeC^/R=(dC1XRB./dV7BS/ZUQEgf_H]E:,?@F180Z
c6Pgc:?,\3,J^IJ,:^OgD8a]ZWMMXC,,WfA1P/W2OUQ;AH=S&)fNfcee7b_L0.-b
D/2ZAN2Gc1[0Mag&7[DVB3NgT>\A9,<3[Sc8P1I\=LcJ?C.U^g0DGWTNZN>e-T,]
U=&M.T\@,HVBU,EA<@Q7&,Y].6=Ca[OC43-N/MW7K@4BZKP4P:VAZEM5LLP6QP36
Ub5;HK-NI)gF#C[#e@(@VV5O81[=G(&TMDZEIS1L7U-6XSHM2AW.EOO]H[CAd#fC
ZgY4GdK1W-EF5cgG9P6BHWV?Q<_=3G[6C(V]U#,WUO84[6V&^H<B0G;73\(Y8+/X
6]#e#O+X-HE^-4JF8[Hc#AXeAR<+UT;c:9M>:I0Z2FaZa/GIXb@&ZB47FB]D<TJD
-JHA92:9SB:N^Lc6I36e2cc/PCf./:UK<X)BOcI7]dYe[R/a.J>UPY?LB)+UJ0EI
A[TO>a&S267GK&@?A5DGH0PO4VXIWEQ=c,-E-N>Y5=(\1Le.T0gS0Kb(O0N?);R+
&0EH;UF1CH+,VT=9ODJ4)EI]\b1L181acI#6?&D;F8MA1@gHdZ?3SRP4)C&_+<BQ
_^&:eQe>e_+f&Y=OHgf0)bG:STSH@KWLeH5FUXKQ71YFfRXKd@JLIEbLOPGJ?@6,
QT5.(b=NL183+g,Vc(]d]MDCKDO4]86(JB46FT=)ZQdN-H:Z6g,73D+\QE<;-+N=
LMT?dF)XM3d:GYL_Y(/a[\OV7J3#830g=Kb-c](E:e,7/cgTfE767(1JN(ERYgPL
Y/Hg<gg:Vf#_aGD>S_bNC&R_OG0#&==/L//<R&?\,e+\M-[;^:F67@FgD]2[P38@
bWS5&V9;5&G)fFQ3W02:aUJ\SS>R4f)/+K@3DNUdb\49dW?0d]SC?==TFL\2N&:T
5+_DB0293]4GWS\)Q7c/([M60G_Q5BFP>#eT^L0TfG@1Vg2TNEb;ZDb?QFPJcT_+
0IWTV2)K>62TTS7TKYIP;>cXGRbPGKUK+):g0Ld):gBISGFW(+L>6G)M_\D^KAL7
\YSIDJ70_LO\26;W(Ig9_F3Vf>Pc0CL+6U^E4<>F^eU<H0PA8ZQYeTffN3<UJK;_
W9683H@bNQ,4W:\X>b,g5C>Y99,[/GcC=-K(gO8V,A27<(.cS4+=D[eX]OEF0SL3
IZ,&H3CW-bdfK-D6=^@c5[5]4=8=H6W49OF,MZJ/(S(/H/5SECV)>>OU3f0??W(:
F<OLZ;)TQWX3&[;bTUB\H]V7R1Q\Y?V463<[HU6<G;SP32_X?V7eL1DHQ?0;:8^-
C^XWVMXb8=M&)ZfAb_@EN-K(A#dA4/g+50#aH6^ZY/5=I+]XBX0[3Ve7>PJD(8K8
23d62?-@,.L0GcKXIXGH;Ub@?H^GeM^/_/b;38]7eEL4__R9/[,a>1c)4^+=H5^F
=\-8KE,We;9^)V9H/cg:U_.K#fB_&U,ZHOc02IL]IXa3W;^\2dW#0K-Ff86Z)KMb
(^S4PV)-UU1FD:;.]<Ie82F4AZRL-b#TTGI?.1eG5WSF8(YU:ab#?R8>/S/)GPfW
:/:COgQ/a7L#fMNJ2_HR+EN[@L^2A>RO^EHMW^Q6WRW8b9gcFX+?@e:f;V.\BA5;
9Q-JEc3VM]T^aCdf\P;G?YeAM5.61d;O.K&6;#6,?c0NRBCUY&H#1EW39Nb[9XN=
\ROGd-/JbR2OGB[3-T:?9)L3^S)F&3U#L>AU\X,/77VCV<^6<NAZ3gYC/L?>2d[[
cAg85>]\:aM+6W,7YDTX-^K9[[ea?;X)7KE^/0_-OT]0bD;6VG6+2)G6a_\T(Ndf
-A4GIL/I2]8+1C-O9Z[T4Fe95?F<.GQOB6-2e6A=71Q:7+XSfcP63KVdPH9a9<:3
=\Z_SIEHNCOcWE.(B1DWdEP#C2Z1dL[AU=VN.3B0UU\(_^&XH\)<O?A9VPU8P?.E
_@CS;YXE>XT@+-MI38M#.EdO\3_;9RV2[+9_GG&\(IVaM&Z=B40UNK98^31>fXcM
IPHW\E7E&>(2^bV7P+B[&e4NeC/.P5&XdLTMB5<Z#@:3JRRCaKC?FNJDQ=dR+D[g
W8=Y090c@M2\K)U59EJWaB3fBU[DNR(QPDY6Z&A?9FUTXW@<DTYNIS_NAK.S2c>b
d?3W3Z&9_g)6OAYE(I@_CE+^W&,LE:)d.A_S[K5RKOG7-JBbNA>];c3f[RM=g)f3
DZN#YH8U5CV&b_HX?3_e@ZU9bROKYQ5YT@=/KBd31UQ/X4<=^IJ03VID]3&V,KT_
NaV^84Z:=_P8bZF<=7[XN)+T?,[Bc0Cf?,,D]4&HW[I43HR@-XeQUSTT[ddLD#=#
^GL8YGJ3-\779PI<[1&CI93bg(1&dE7VEN\T.e6G7EL5Dee:DT<63001/Q=9e04c
>;??ZL221fV;B>e+Y-S_F_aDdW>L65H\4d.N2eDPNa-RXO7SNL&]?=CZGf-=+4^U
fGRDaG)3Eb9HWV@6D9a7):>RB,Ned05:;eUQG(76:,)N/2(#:])Qc#QD3>fYL<^Z
fB58LMGF+SFF=aC\I6([/&DOP6g9Y3,&IR46L[dR<=eg@4^5EP?XIJ97J6S6FQg[
JKb71UZ]faNW3T?d#W)AETfTL?g?#>&Q(F3:.ILd7BNdZ96M+P#^0YY>9<9B[QH#
<^XbG>[fK[/FVd=\+90J4O5>IN=J)LC)NI)C^8T32T,YF5.Z_2W9A5ZZAecYeV.A
FGU40PLF;4A]d0b.?aZR]I0fME>dP5<[K4:?d<&OBf/6-@T<cN(DfM1#9cLb(eY4
fHNERg[/a+HD=(bGY-I2.7ID9G1TP,L,F+?^^PNZDP9(L\:C8SS./[P(-.-44Y,]
AEO]+:P.SJHc_HRZ9-e(R@E7+Q_2b+CC;1-;U03<JdR6Fe(^8FcPa+6QJ9Fe;aFL
@6>ebI/116N/XN^T,>P#0gZaD0RUfUcD_f+Y7LS8#J7B?SK5HO2Q+?9ZIQQ62FW\
K9L^&8>d\;;SRc-;OS^V6cS/81\A;<&;8S)._F80=>#35dgB->_:EN6aTXXbabG<
-UO_DYT?e4?bPQ9>F4C4DJTMf>[FTLe.N222UI_U1[PM1;#gSK#9F\B1WGbS:_?[
CZS_U0ScTbI,EH8Dd74a&W?&:W=DR1U4J?(81UI8aJPTX7]5Ig?#HQ/b7.dGS-\+
gD3L0[SSP/:A1+)H/)#4]aR1EV4.,Z(Wg/+8\+0MXTF^T(])V?S1e1DJ1;J93a#T
XYI(0SQ-])_gfJC++A@2SZJ>9/OG<&SFXOX\6+7L-V@&4U#-Z8DSG[]IIc5gd)bZ
<5d;3N86AVE(J8.C&f,?7#D-aZ9J,P5B/Y)+EK:K7g4[+^9B#P=L>^c#OLI?D3(=
))6UP4_+EB\X/;cQ99<(:31J4+\S8P[VTAB\a_I^C3<Gb,Gf4DXK:V528B\W[APG
CY5YV/S-bGQ6K-CXJXR1F+1g;;ZZ7.e0DO9MV<Zd;=-EK#CCP9+HNf.PHEd:W0XW
JF)5Ef6^ECfF#87>UX/f)=,+aX7+4/eUTX,E/K4&)AEc4Xg=B/EQF,N5J,1,[-P8
QW^0I4[7O&FdY_=_dDP\DKKTY9g+4[1[VQ\dZ_P+455>fT6A;@/Y49U;ebMRf):(
8,T(a6)17MV+dOQM\+P69./:,L(>B<-@(KSNA52;@a@eU(:D3;La0^SdSBSHO.Z4
&Ae_A26M=#a:HW_/#b1YaPJZ/a]V6fD:]F+@_B:OA3JR@GB;?7eeY.Z-:Y;KY1Ag
PJVDgJ9W4F#R\Ad,^SYY23G#=C^c]]DQVVJ)NDKg,KC#;3Ig0^G;1)1Xd^XYTI:B
)3PLYbZN1SE=-aYe9==@\fZI7+-dYRH9:<8BXfd&B35)MBFT3\7dQ&9OgO?CMSd3
<<\(SdQQS5)BVH?O(7,LGEV6I4NgH+6/]g</_B[c,TaD+Va^_M3c644)VfC3#WU3
b4+2H@dNbV4KM)EFPC<^g<bD.UYK4O_\/3:(_c7SLJdYLN\<[K/FFK)(/9B&-V@L
RMY2dGdRO,NP3NS>&dL?0(ZVgYZV(bF;C<4\6K(6G7W];2fFR/GT3#&e,.Sc<Qe?
Ea]g9K47LW4IE;F+(--&W08VD<R(9KC>3@/eA[>1T@,ORb1+SL=6+J7VTb6+J:R^
(E)@QW_Z+@<NDK7f1ZcbH6Zdg9Z1DE<DD.D+G[J\G:@J-G,0047ZB@6aZI4?A&67
]<Z^e(Pb^g#&fL\9>7C,,O8c\1MgT8b#_MD^>_1S;J?(6Q-1Tc33-X1&6A?.7Q(V
_Q-2#QeTD=LZ.e_bV)Wag2^bFNDb3bHbg7_6;aW<)U^2.b@85)=I?T@UfV/N=5U9
\GE6DWII.e5eeg?YM-X0<K9#J/)2EX=-J:Xe97(KT.@Ba^a/D9]/,A@^>9&L#&^>
dA#JD_R7f([Td4(DL43V.+XWG<GL6TL#94@<EM;;[+R&;Nf5B?^bUb>/HL.f9NG8
[M&)(.g,\O=9c;NTIUfD-[(gV?GgK6(<76:?KF#,>T^U15+\A9b2E:D1AL>A@b>7
8eT+2<JbcZec)J(X2;MZ)DA-SN>/,a7P#V@>127cW?a=KL<CE)HB[5H]MfST9S)a
X7CQ7CQPYcO]CMNBNE9d_U=-W(.GF&4[:TFI1QZJ6JF3PDU7,\8AF?4=]e^)M#<b
?:]_9,J+9NWN@g?bZ+F<SBX>^SH.N)c2&01YZ83RJ#BV8ZJ\DJ.BRD6I\\/Jg+A]
e@c4dDM5gNV7PX7.eM:@Ff3I,H;72[b)&,a8_@G#V&)1YV0@@Qg6A>BWR/D8/;F,
fLLYaa[WO=g.gC[V1Y(::K;G+U91.B)#+:DS\BX@^[6MdAY&&\PQ:C.QWW_P(,J[
NIXd&+dXf7Z^BFSNNVc1/)9R6e.QG-\8CL7/[^^[e,)-JQ2]M^,>KO.UaYP2YY7d
-.,J+Q&[R4c-@bPC420,S\7-+_SY>)S):V+B[C-Z3K\(2;?Taf-\=D/GJT]0]BKa
aY[#JdS@#K3\2NC>6bf<;gXZN1&aN&4\2eZ=33&WLK2HLEaa.+R-8\Z]fadXc39P
2RF:e:S\c47b,AaXPX5:?+T+RO?;/I^JJ7c90Fb0S38@4(QO<3/OQXQ8K=9G-)])
#/-?BTV_OM=(3_?:LJ7@:((+:M+;@)M/.::22]bGK,GecZ:ZeXI/a[1PH&#^4[b_
S(&ZHGBc<C<Ec[8F]BJ,Q<SJ_CZC?=L=6#4#@;K=JaZBX=@A#RNfY]\,(\Kb<Vc.
3Q?A98+;Rd..X?ZUMdX8.(Q2L>=d#aNO;daZKZT#32(N:X]CU_,g1QC17;e]55,E
LJI+6FELFQF)79TX66[E_A=PI[X509W+X+]f-BT5TbK-,(-bZWgf)PCJ:?dXDB=I
ENS-cAY4R9N/[?=YXPf1CX/_aV1[gBaZ2E/fWVQ^0d&:1=_T8Z8;B)>N-:a;F_+4
b(1KSC1fe9]5#c01#6061cY+CS2#3SOO+8eR&e(LVQ=<?8TfB)/]J0D3\GIDZT2a
&^0[K#(GN&>Q&])2H?E=D&6BV-)IHHO1&P[/HND:;BXc6OW5/-7<+0:[2_I&Z@W8
:5[ZT5E]M/fV-T-Q)&g6@d7)3+MOSbGP?_3Ud@5AcLD(0_7F6EZ1G.20HKCB_O((
(ZX9/fSMa4dUfaF]__:8-A2MYCAg0Y9#93Cde\L64H<O#W?ZbNZ5:AgMaKIG,?YY
fBFW.^T31;<Kbc;;),:<W3H3-DBM&NBWfIe:e/CeGV+Y?+FP)#SOOPW)gSUPgHeb
X),(LBf6A.[-7.LCP-HCVIYQ@1VSEFT]OVR@:g)R3US10R.Ic]?I[]1]ec:b6J,F
T(,9.(.@\7D@)L9QDMG7gIgL?HU@EO_ZJI)?[TL/<AU^2D[(g#aH^4J<4Te)D>b-
dCV#<90ZF[>deP<9;^S,a-Z-_R03UcUd=d>N1AWZJ>)ZM#U-BAQX5#O4GLfS2&7P
a9dR##C&?NLQ=O)e\4,+VGf]:\(gFJMeWLMf<]4(Va]1@@G1]K2H,Ng4-9fTE-M&
^0:J;&9EQZRH_??]/MK-fML/2S)a2W.Xad<Ea-V8U0(<YX2>Ec<AA=LgZOH2QS55
5Z5D/1[\Pac:MR4MT&SJgCaa([&TY3Acg?WYVT=8;];)I(M\XE.E7@&#_YT>@&(S
U7L-0.S/B[)F4Q[I_gU+S=Qb,fR((G=02;D)9?62e+L2J0?)-,1cLcWIAKGQd(E]
3=0_..5J<f;3S.E-a,:&fKS0RS-SZE],/=N?/f9TO:/&F;-SQ&bV4&5#54L0XEH9
a\Rf+JXe.MS31bIDWaVcXXL+0>:^T23B#CfXc#fW1O?D>>:?ga=P/OJVLWS4R/9T
;JQ.1OcKLaRb5N<cL>G26AY0]OcRP>[R#d8WEEe+0Ic23.,e,)0SL;?5^TCC2_Vg
0CNU&6Y7Q#b&UJI#JZLTMDDNC7B.7eLg@V#O65,0+L+/[6U3RSHOf)5\W+Rf5L^d
:N=;6HOI3GUP5ace_J,f^WBB(<KKPU--GG_7GX5\:YU8D3JFV(<3a13.d.7EQ3QA
6d0,4>^87b@WfXVG->S&^,2d2fKS?K,JV=(#VX<+/Bf3-]X#2V>#2JbP:-)G>U6+
Ea_=+V.B?7R+.7J,U@)LRGB_bc.-9LZg=N8[,-baPP::W?@YCOD3/[=bR<B/eg6+
H.TGfg0:M<?adgfRL-[K??M,M\[g7/@DBQPYVfR.a)@:9[e@CDT&NBH4+KG?&?=9
US?=^B[S+K0?R&e?/.3=,\RS0>=bY/\P\6X2IGV?XV[YY?)EY7.EK.>:<;D)-KK.
e/Lb2Ucg59dN\@0OLd<7[]<8GHdI1P^2>K>KO61G-cADg[bK66g9@CeY2CFU8bNG
]-N7<\2]ZZ66b?EYA-a#&,HGWSK:16O#E>-E)HDCZ(]&.DU+=RR8.)Cf&9YgJ:dY
@ed>1@2f&;R8/?(5^F8&2Q1C1,I7]SfZ32AYVcG2S:/1,,f2).\.^SBYKa+HAU81
e<\0VY_.V4BW3HEO#ZRS]X.;[QX@UA3;84I[_2,T19D?g#\7B[.0//&8+1@4g+SO
=g5FA7SZRL2dKdSE]^C>2P[,O#FR&bdI#0IPVRT,B:JW[+JWU2JIE30NL(\b^/Z0
]8<#B+XCCM:\W/SNQS)1?B3CFF1=(N5DaFCL,,6VX5#371QFUH3+P&ETL[&64_5O
Y[7CK?Y:JOb#KD4P0_d=0XGNb@5?LGYIGJ--2@;TRXH?TENYfBY.Z)Q6ea)&g0UI
52+;JQR2VeUUA.O-I)0K1b:=5]WD#Mc/7A4#Z9B8R,UA70;&K&#5@d;8CK6IFcHb
d7Ea/:G&=E2TTUc1Je5MS:#[QIY/eC04a##d>6UKIV:F=BCW_X5eSE7&8V57NZC=
D5<;8gNK?98@67OZF]^=WeJ.[3/2[J1\9Xg,T<#f1\G0KJ[b2S=#(V;Cb0<K3TC,
DXEf.fdQ#<-/F?&9LZff:dHN1R7LZ.EA<Xc[X+V-8Z@BDLTT75e^XAUQ7YJ3T+?U
&eaL]bgYJ0+(]KW\VR,Fg/,W>MXN,-RK&=RY^U[XGAaE@g;7^Sa5/bXQb^1JU.GR
@DG8_O5[2=IU(dV#[(L&=Q(E2R8^:PeAcWOATQ]J:\3PNXUDS/]Da6fHU@_cD[A?
c9P:XI\#eUTM[>_0N=+3dI8Sd(HgT[a6/4_K6?,Q1^]^:=>WY/Z6:E/_VLO>^>GX
dc6JcMJ,?PD,XbH/f,W0^VFZ61+MMP^8BbZ9,02F9ea+#,UdI/b\c[,e-fYFBSH:
Dc7&[5Q=-Vf,SS)CST&ZFU(09b]WL.>PJW8KFOf^X2Y1,QCS]EXb)fPI@<&V06^b
FO>WF=7V73T9&Ud7N:5Y#Y1d<)Uc1Y_KTQgT\Wd\FX4GAPW^3\NbBY<=,F>aXG81
07NQRD1(-a<TJ_IP9E<#\P.Kf74a[W?ae8F0@>3)XP,??[B(42Fg+Mg]LM@[5]X,
].FAMZ55Ue:d?RL)#B2UI=4(E.dK<1O8D/0RFN74W^CY7F;GZV(+e11CdAV4#]57
R:1-<(?=IGRa:Ng,\HN6X4V:4UC,?;4X>Q]23E@.IOT\OdELXe<7P4LJOZ:3WZ9,
(Kc;?&CD&6<@aTefT5S^(SH=&@#?59Ug;=;Z_RXVC3R/&9AY1FT(C2b,;8C=41D2
GG4196SN2Nd)WfY1XfTOLML>LaDA55\FN.<\+W.;Ag\>3;6Ne^PK&RW2fJ6T8;R;
Q-H)QdW=4K,0AQCALa+XPX7[;)^Ic^QSc?\V=1VQ^3\]b\0E57>4,e_7Xf@+2)E4
dK3-2?0^e]Oc7>2FP@[1Z0V&MN@QEQ:d==ee#+:TQ7&GOV&GF]IGI+AUVD\]KEZZ
O0OXUO9@g0GSE)?&>AFOb/0X4J5ccB6@OQLb6235>2U\4GY27>X9f6Ie\+S8&X5B
98FU,&VUBKeZ-GES&FaaV-b+Q?1:4_^OI-1];DFeWCUUDX1\EEW/Gag2<EE_a&8a
]@76HF4_?T_cg6;T).HA6gZ+C=#><(BP3[L.^;M_13R.?([(..,;[Y8:eA\&L,KM
F2.Z^ZFTa5X6HcKa.HPLa,6Bf/+Cd=UE6>B=I-(f1P)8@fL?dPU?NE>SA5W83HgM
=\aBOOUUPeGT8@?5La0ZZ\V\1M:A9;U_^1:A+b(Rd[JF&eXB);O:79Bg?6DDW8;_
g[F9M?72FXGeABAEDTc<eNT&B=eX>.FGZ4,]>(M8UNf3Dd&d5;@\EaPC./)0gUcd
eYHcEMg53Ff;D=NP4>Ye./>@K^7DaU,HK&M<\T:/gO\-H6d]DU[R,ZF;f)^,8?DU
&6UBB81&00F1]V&P:TYea>M=G@<5R1]aTM2,)4dgG_1:U6E52RH7LWH+K^4Se26A
;agDUZTM0F&@[5B)e:/Ccb_>,\f:6Q>6-:/M?HEI/F#PZ04_W;V(FeL[8Nb/VNND
/gV_;IdJcTeH-HJ-.<LRSbcB,c@SWL[)GP+9La,A-2W)+>Q;,HfW&9;5J.N;R.J(
V5P41YF@K,KD2-cX9abCNf/+Q6c7G)ENPA(F-\;HNZ5J&#=H=?@H]KeYc6)V:&Sb
Ab.TVUcS0f:O.5L2OR/G0FAT>>JP(@\K_R53>=+U2AEX.PL@T9Ka?@[V6K@)&4/@
9<CW;7GJ[Q]UBSPDHXZ5a<M^9^c=(GSYU+d#>TV6JeAC&.E>](gY>;C(ZXXb^QF,
E0@dU4XS<H-FI@S[D_VReB:ULT3T4=4F#SIeOGRe;;\]RTQ<()J?FBEWEJfR#NDW
EM&31#dVY9cPUW\cWSdPQCYX@M=LSR9S)GF\ZC=DC]NME:/]X9eK,a[\7Eb[f_NT
WJ^4K&M]IbP?[3aB48>#dK]SN7/K]g8Q>_64+(E8ZWVR?0Z-4,,+[ITZ/DB2+0.T
N]_C_AXJGLEA[G0OMS/J1Afb\f21;M@))Y6JT&[CL,VXXC<^&4+U;J/C@=_EHNT-
3S+;9&fTK,76gS8U-;LY4Q<ce3<C9b-2KG?3QM(Z@2;QC5:ISR#]U@[EVU<:[9)\
Bf>/.GELOP,+CP\BO>1#g,W-@D#6892F.>[<S,NUF>^gN#(E@7gN:#KCAHJ]T\&A
g8)5Qb&WG&VUXd9]@/:#4.f-g5<RcLVgTc_RT@5/f:4G;_\bA#HJ_GZL<KeDda7e
0Sb.E_M-Y#X3FHg+=J=413..F[N\ZO7bgXR:-VFN1Q_V(U,f1UYUa/6bD7[NJ&^)
>X]gP694.RSTVf<[/C9ff3+Q-T)/@2[CPFZAD18?.EADN0WKC7YS/KBO@5)-369>
F)0LZCOD:)OV;aLS:0ZL\9DD@;X\0R#U?_PA]F+Ug=;cT;>^d59eR[;Y?WYLR36;
fa&VKC6cQ/A&.X07D]gH^(#W7)9UIg+[?<.WNf5/50=,Z,&NfBVE4VYLGHH[9=dL
)LY4YH3JNc@\+?9EgJffSP)0&deAS89gc_-cT5HQVMDD&c>1O9O&6S[\Sb[?0Za?
ReQA:9,c@&Y=EDO-<E;_K8\Z/eCTP?f-7,X25Q&d[&g/BH_9c/5e,^SZTY#2)J&O
#RL-gTDa(0),-R>cZgX7<Vg>bBT42U;Y=GE=>gUFb0(?)JZdXb]?XDD20B\N]&4a
aYbXaD>ec2K=gI)M193gJ8;9/8\/F5K\P.D>c8((79?.24&Vd(4cJ/7:,P+a;I]G
<(.Y1\D3bZTIUA3#^_[AI^VL5/XT#QOJTIc_6]-b86-8#<>/6\)R5J+V9[VGdX3Q
H&\3U,H_#AQ9Q0]BF=EZ1\ba]+gL2.Q9#6]HFGbVLeXO.)0S&(:UaWF8G<(KYVHS
]/0<b.M@V(a?[c<:<O[DR2;?9]Hd@Kg38gMX&Vf.bS>[<[BXU1Q]X@b>8]()H.[Y
2Og;FLH)cNM5DUYX6]e3eYBI^M6>g.D(fD0Q?f,=E7BW#Oc/;_eJ2f6<A8A(]8A2
OT.5fA=<2f7UF_;W09+R7\<ZSLBLR^L/f:D45A2A8R_DOZdO/feT&E.E;IXG8_=(
&0bf->];-,VB+X6V>W?<<886->?W?L)+HE#.T_FFYCL.JD2-fWNEIL,J^-3Q(ZM3
E9FW&1Z<W=bQ9H?>L&>YL-9&X06(Q@8aTB&P)+&PMTJ^_G+=L5dJJRS:?)_&D[M/
>6b@MQSHYQPC)S3?L#2.B?S=c_O]]B-B)_Ud?RSN\Ue&dCOP^e(6HTL=&80cO4fC
J<U#BJTCBaYZ<J#5XOK/]R^H5:RIER3a-M)]K+gN>g-VRd2IESLQ8DA:)H(?/L43
A2]WWLSD/e,gD@EPP[T5:^e-+,L:[:=ES1>U:(E?6g9Q><P&H@X//E.-S3?.,IB6
;(\BU9JR555:QAX57fYK_WJ_>021[-9ZF0E[GA?,\[?GD290a6BN8_NgNIf)&eK)
,V;>79413c2E9QK\I>YTBE?SB&=:J,eZ@B:&a/7/RN1\##P:DT.M99BT;6JNX/(f
6_[,,;AKfK&JXTc2@+c^d8>LPTb0;aGFDQ8aYBf]TRLGSE2^2V;Z<>,?D@<6WP&Y
EB=-a/;SJ_W8JZYg[[M.Af9GEWUL:VZ=L5WC9cdFC(;#YC2=PRgS>XeEOf=>.ME/
;8\9AgEbB?ga+PC&(#9R\M=]IcOVO)#/CO]<4C&D:3e0=A()529Z9([f2RK>GQ5U
OA52S-5dEfO?=^bg3THBF;1e3\<:+INg3U1-0<,W=(7_?;W<R.(^/f8XU+;Y;B,X
O>KLD@b\C1I>7SETdf0,7C>B9M3gV;g5_Hafd?J1:M/R)2B.FN3;0PDWDDaQQ:H9
)>>O7IX8@&ebM;;]79gg?a-5=>/H);\Na14JDOGe6Q/43^ZEe-e=g20]))B#SQD;
EKaQ,de=eFZ\bS+3#QJM66@/_[YGDFC1UYd<GN]bf&9JDC8S6M,M/CS3&fK9;gN^
H6&_+AeOE79?fH1^eg]1Ed5JI,1aM,WQ2&O10:,CZY)<49P.)Y^JE^dTa;=7Ca-/
#8;)].2[:Hda_V4[&=NNQUZLH(I\8&c>,?Z1U9VeUJf[;>M1=/);;T#SA4(&/L#O
_\>MUKMM7-bcG##9GDLY3f/(V4QNY]3eBXNeW1+=11^O7dFG9^MT/:AOdP=AWOCP
EGJ+)0>RR1GKfeJD#;;WPd4=VGT9.3876]N@&eFQg@4LM3\+-91e@g8-/N7B^Y4G
V9UC=A_>ZU\bRe-KTG_KA6/@XED+^dR4&S2,eb&38A3W<a^2(g)@O?0)@AMXZ;F&
U1eU_7L9Z&bgf;fE=8+5SeUf1_H0fBX;;XGBQ-d<8^@LDK[>F<3N+CXf_6e2O=O0
;I/4.H[2PG^]@@^c)5201;&fQfSY3)RdWaS;8dEd6-5)_6JHW=8NGd\:=dT0CQ5;
#4?TL\bg.EE@KZ)PHC86O,#F\YR<Y^Icd9+<2JX<f>1f?[)=0G,O#AT9MEPZ.]\.
RWB&;P6HHZ8Fcg@R;0TXG,&UT96#7AQ<e<KP23V@W^]JHXC#1T[SRI=K95VT&V/[
YIPVe4cAB@G8RELdad]2/-@N,TWH^<;NG\Za9NHA5@0>fR3#VeSZ>[,&aWc1N+AW
2JZ8a5X^DOD\[HI3Q5IRXg/IQ_?,a+_4NI4@7@+B[5K6dE0E5bYEY5UY6#23&>B=
1-6QH5IXPUeMJOd:7)TL6+Ge,\H40&X<8;+>G7b6=L_QZTMWY9.J6K8A5UFY[9ce
[H3N/;AATe&=EFQH8HQHMXXAMLNT&^R-5+O74#Y;;eV7?,0BgcAdQ(Y)\g.a3GS9
Y>c==d8DIRg=3J4F6:6#?R#51]HL4W[]V3MBL,TVQaA8b@2Pd[g:4\:\[@QKb8DM
(9eOTXV5FU5?1-e7>,:aG9DM,H^]7N:NLE&0LB(.a6Hg9<0&6c8UJF/ERE0<V9AU
PKO8G@(D2g,46.)2c_8^4JfD)K:LbAgPF1T?<3#?/_?R3dg0R:f\Ud45EA(Y@<3L
FH2]=)ZfQ[Z624]D^_F>d;5LFJ_)6f,V#e+GUN)SA?2T[UAN4XM0ZZ51/==6fObZ
gdU?.=BadEa:M^M7A-(\NU(e4LL;H-Kd8GdLWL2=0([5>[G&]6T^0#EA5^@g/c^8
F.<8^R7CV0\T?XT:^G:X,RMGSLS0KV1)8fY=NgM_gV?LBcE/>M0^FWeQ/<-Y#-6c
M<bGQR[(]7d@31R5dZ<AL8[N-AWM/24VRMO1UJAX6X7#FH[M82>>^>Y4^J<0D6Z<
[T9-K,-VVVN2W2J)3?IPVQ4?&IYC7b1c;c(^/O+T+]TdKX1?N)4;6R@K522P+CU2
SVR5R/=Dea_=OGI3G^DD2M4,NSWXF8eA=Dc)P]=57Y_IGfbJQ,CbP^&dADOTSFJ>
?8Nb,:,&VSMS+R?[_<,R9RcHP=U)UL[YEU(CFG1=<.Ad<eNR\R#.a_-Y.WcN,93J
NRZ^8PDUM8MY,E\,+UH_8Hc2/c;aD61\JU[6>U[gFg=F\#:@B3E@&(,].HJ30(\6
:979eNHFLA.?\/Y9eCaR/T[?KNH4#/L>f(S^ZS)DZaT]4S,?Hc:1YF>5e..).O2L
?=2;?Ng-2W/@TZR?0bA5-1<ZAV/.9^BM7:L8A(>LJca9=]UTKaN70/adKL]A.LRN
.691WU:LBNI(7#K#XKX@GPJ5V+.2_:_beMGYL6(2WA#^U1#?4U:Dbc+/7_PT\X&=
7@a7,Z)f5WC/X5G,>Q&UX27,g5,a)Qg#.R</5PccX&1\SWX])FU7Ag7N/ITB>]V8
+AG;_IR[A)LJX?I7<?He3eQ(ffH^bAe#aTMf>QPK4D_12D:K=a#^GcRD_<cObRgf
68;2g9d=FJ6,JSP5M;5[GaOX0WLYaBIQbbCIN-X4VO03L3.=TMdF21<#cOG>?[6;
._,SAS^X(g+C;LSg1V?bTCHL^3<G<_ZQUIN-2REL;@cP(N4.T@JNP-W2511Mf]RM
S1_fBSG_Y6&:HG[Pe.1EX(@b7<4OU>BT)M@bc[ETVC69;Edd1OOB^E3WD5HLGG5P
R(4,N=/:IVET?+a#4]IGU3Ce:0d,AV#/\U,+B)M?8T7=BgeXgZda<R)a7_8IKEf[
ZbaVFDc]A@]aR:+II/(Q0PPL6F?)3M0>[;.Ra_(gd)>IQN[O:\+;gGW5U:e]?g;Y
?/8VM1Q\BB27B2gH)>X#?dF#&SWG5SZ.VDTYIU4YBVW6D8GPLA(g7K78;:)4AHf>
ad4HJcgV>RS@4KbC#MJXf/0?dD50X_\N,^@QI2)GLKH,MS2XEgB[Z0\::1\IS,YI
<M=3]YBLDTCSMNfL6:aeG=aHX39:G2:RNdeWOC-+3)LDAeCPe-<3b&D13cEg7b<a
;6-:Ud-T-)2UEQER&50M(XUE0\5J8J/P4+a7&GAXU)?)@8=L/Re4/-)b-\^f7=[#
;.VY2b4[82Jc)e;LZP<e@2C>]L?Yb]NQH1C(b<9VW?0B6,ONZ<@HH;)F#SU6A8YM
ZSD,3#[fI71?APWH2]7G?C56DEZ,LEad9,=&XRJf#1bL/334N[=W9-=2=6VL,3(D
2Zf1?L<Z\U+1T)@&eOefEGe\[=a1D^CK2X[095#86;c_-=1d9bJL:O.aRGT0(]E5
9R6D6-e>-I)gMdd_M&RAR5MbI+)(2KB.U^c^>U79]B4K<(1S4<C4OB=e,1c4#W(V
YSGG@:UgERC-/W2O<J/6P/^ESeC0PU_K;LNce,?GH+_e4V5PG32FKNH_fceY_dA@
8WbKE[gD#J.MJMH8dW9\#RSec0TCX=FC\gJIC;3&M70.cG9(aP)TReD1gd8JA)JX
TG]^A[N6;PB0W\f1#-553@HM;=8g<TCCM>P2/B<J;>UaD3I@_4OBg/:OeZe?<HG.
b\_]SU[e=V-B52K4,JDS0b)\WG,9,.Wg5Z(Z<TO,[7Q,NEZ=7^aea]Q;Q_]c&_EM
FTaT(#.N)&9/)^+.Abb.05M0GL<.B&1?5+dKd;SMc\dbLEA2S-Zg8)c=]I9\2aRf
+8BX^WLOKKZ06gALaB+4gB_9>DRVKOK;L;0H1+3XXX5PM1aJ.XDBR0CCQ?.cGafb
7<_<+EdU5?I15&;SH]R>dg.K[ME#U],HfgK)b,THb[YT71_K_NG-X[)4C?R>UZGP
]I;b-7YRS:Z8.MOVFC9RQ48VDFW-Kc5IYd4:)3S/<42HL#[aD#._:Y,:b9M?IVSJ
8A9V[caOfQP9DL2E6<VG49ICf:b<XeF.J0gXVc^:3;M0a3OJeC5f3IcIU^6<FJKd
\\56=C^a6LM>C?5NONbZE6BN+:b95F>5K#cL)O:4YQ:G#Z=U>07R7MX[;29.++2\
OF;ES5YCc<?S3,07fI/FW\Xef-\AI.be)b8BGYF\\_^K8HFVKPIK,2FS[NHe/M_E
MWUbX=/?EH#B3.9(JUaNg(@BCF^.F?FJf.3eX][3F<_G)g[/X\KY^T3J484(+@@O
04DTKgZ02S&7Wg3HbY@U3<&^JHcD1,2Y7UeK:AP3bOfK72OW(]Y3]b\-]/[0242\
^B,\(770<C(PaDPIISL00S5.P=&WX3f11/U@9b6_fMC#+Hg\<HW@d[[4g#<KE4TT
SceNI;AN+(Q5#>\VTf@NE<Q8=]O_QRYa4N38b4Y2A2UUc4//fTeB;/J0/aHE^eEH
Tf830g[-P>f&5_HHJKS^R05gIQJMR@2ZZ;/RDe\/D1(8AW]OR][Z3#=fE6H_c)DD
6?(0VJW1QIK)^./J?EQbV,O@Z0ZN)B6Y@C#/JZ8DS_5?<OT5L#86)5SR>Jfga[E^
)V<@L>FbBgcg,-Y)fI-<5?DD<B-8=H3ea+;E7FZbM,PI)I\S<)A9E[Ke6RCL64cV
1_D0G=,0C7QJAaN\.FdL6Q:E(Sg(A=B+22g3Ecd\f#V9A03NNQZRV[E@QG3gd/L,
=Ne-ZWLT-8^g2(Dc_Ie7[S12f?0M6?:f)1SdO9YP+_PReb81Q=RPJTQMMM7H05JH
_C_WK]HfCdS=E^,/E#]PB:.W3V[_[VHa44@a7+Qd>N]91?agMCE2-1CJ^B;(dHXc
.U&b@S=Hc@&J9T:(a]RNLKS3+W)/DTAZ4P4DJ9b;-S^W<&b;FV(<I,MJ6LdX/TQI
7-VO<Y.JI_T\AFTO37&V0R#e3;2cSXVFR//Q=D>?]\<MYZKSSQL;E;JeGL?O.,6;
T&^L8)g_+;)<<SeLW4JS\\9W7fG1aZX+_[J/@-SY,Cd_X<T+Ad\TMJ17,,Q;-_\0
XEPJN#bU81GTN3Y8Gd\UdAJDb[RgHE\;D,DO<2>ZY,)cgT4C8WM;^]bK+d5:0L,B
M,V;[<U(BY<(.41E2UUD#ZW,@D&<E@\=g:eNB?LTS,/b>.NS]:U(V<B=J>2(;^G4
CL(?&6H:\eIM]C2J/[JC=LO>@?dPd-Eb4c[F?XDgZGeb+[#,C,b3U(IOU)W_0g,[
[9K&4.>&M6VO0#gD?\)Z?-\UEa[]4:b(>(JbR/^#MY77MeIBZQQN[eGKf?b.d4TV
G=>\P465/7Q=R&cWgCO[KWYc>/^?)#FHN?f-(\<-f2(PV#V&(.b)#.FQ>#aL92e&
,Le2OMS4+a0OYab.TCJO@871XX7BWc^<0]4IHDR1e#H[bD8^D<F<aW#,EU3O_D>^
=Hd4Eb5-^/#Nd1;b\b,8K9X7/T./_f3?IgJB^X8KY-_PWIKIb[C^#:6V[&H)ZVd<
A27&9)5DH#/+&^GB[K(RPE-T,93:fIN7F9ePIW+6^3c\(O0e#.:5d5EMF<V2>beA
=:LO0X0cXE1O99f43NGI5@XX#D]K6/JY.fQG#&V,Z?/9@F#S&:()ND)eOaSa8MOJ
<(9>I<b(1T6gLIC5JaY:9)V,=QN;>G5T-DJ?bKQNS]QCD1JH,+<b5:\@.GEX#aD-
cCT(JcH2?Wg66]95VZW5NI,W&B,JT)^<4X/#B7:E(B;KBOQb2T5H[Xb\X>4/(M@G
=:EU]F_C)dGVI(Q>2H)WVac8U0)8XWPEHe[)b)H)Hb5b+HXf&]996:^2bHPd&Z_9
#0FWW.>8DT1UI1SPf6BC5GJ3d8._d78BC4R&2)JL3JC9)-4EFY)XO4,BZf;+>g6-
JJB?bI6aWA+d>R.IQCG3cU\Y8/:W6f@]8<[Gd+07THE@+9Q#fKde9M3<9c8Md#P-
J]6L6)<DT<F1<@6C2b)c,>PHUfZ^I)eR5I_a[,@c2S]bOaN^RQg@fL0bG-_&e;5c
2(]RP(Tg&.SLY3H5TIN/5bf+6Se0dfgXZ0AJfUg@-O(&9J7F6<7ZC[-.3MZ)D28b
&0(<#5(^6LQ(YZS26=:b/97G.;:bY6W@:LcREf?5.F_eGAE:;d6?P3gaCW:M1c#O
]59NfMEXRAMd@_<H;3B[\/VEYFR]PO\/]#YGN<Gb\C546PNN5WTB^K,E=9_TE[OI
fAaYfAJ<_d].Q\>SV:f&/:_b-NX[Xe_^F9ZH:DX)?ZW:1Ib,Q#12^4>K3+@fZ26(
9F[<WA&L]MSS9]AaT^:4(]JBW7BWRe5X)>2[;PCR\bRY2KSI?#LGbgd.^1]D@2YY
6X_S_.g.F?40fWfEN@QV#_[,a=&MN/dQ&>F[:=SI0H4Lg>TN^f:H5@9NOV]>BP;5
5>F:Jb&a/E&Af(Y[eN8e4-J8WDCV[JDWUGE?<_C)5.[.22JQ)Q<Ib##/QQfBd==W
Aa[D4KF3O+O6^HB62IJWSR?-f^:f(XJ0Of30>IfQU?FV.[eTcFYS3Q5UUB6@8F20
&)b^@bMc^P9Pa;38NTR?LM9[PV+BH2_G-9ffBHW>ZBb]I>(=@H>-9J++\U]f/&Gc
75>-N_RS]WQ\/:22gHJXQ7+Xcb7KZO35EF.K@=fAMQ4MDT8<DI,C&?;CT._[X=1+
>_TW0XaMFNGS(K^=U9APR8d->PQ^HFZPAEHJ1#g5PE&-LA;8Afe_?PTSAZXVdD(6
+1BJ.>@0XS(G?ZQJ(f:fdSI[?</_SU[bgPH1,OUQMe1FX@XF5<;gcZT)Q?EZ^]Y/
]6=cN:aX-N^=-ZD3DKG&,0EE6QFU3YI7+NeFBNNb;.CT(WP,)<D@B4:OV(-;&e<g
3_.<TdN^[N\S[0:FT-2__FM<J<C).daU[34eeAOd@UDf3C[3>D_M&fOMf^Zeb&DT
8RYZb4Z]U9bZ/1/)@(5/.Z(/5,EGK&)a&@2V#X-EDB-^Q^K.[825G[G:W7P&//2N
AE6>-4[.5-g:WGDX24]RF<27gJ@f1Ug\HTARXR:A8HbRKURUPL&H9#3Z2c@:UfK<
1/fND:L7]CS:*$
`endprotected
