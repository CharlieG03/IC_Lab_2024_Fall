`ifdef SAMPLE
  `define LAT_MAX 10
  `define LAT_MIN 1
`elsif FUNC
  `define LAT_MAX 10
  `define LAT_MIN 1
`elsif PERF
  `define LAT_MAX 500
  `define LAT_MIN 300
`endif

// Modify your "d_DRAM_p_r" in this directory path to initialized DRAM Value
// Modify d_DRAM_R_LAT           for Initial Read Data Latency, 
//        d_DRAM_W_LAT           for Initial Write Data Latency
//        d_RANDOM_R_LAT           for 1: Random Read Data Latency 0: DRAM_R_LAT Read Data Latency
`ifdef D1
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram1.dat"
`elsif D2
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram2.dat"
`elsif D3
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram3.dat"
`elsif D4
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram4.dat"
`elsif D5
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram5.dat"
`elsif D6
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram6.dat"
`elsif D7
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram7.dat"
`elsif D8
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram8.dat"
`elsif D9
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram9.dat"
`else
  `define d_DRAM_p_r "../00_TESTBED/DRAM/dram0.dat"
`endif

`define d_DRAM_R_LAT 200
`define d_DRAM_W_LAT 1
`define d_RANDOM_R_LAT 1

/* Dont Modify! */
`define DEF_OKAY 2'b00
`define DEF_INCR 2'b01
/*							*/

module pseudo_DRAM#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=128) (
// Global Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [7:0]             awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [7:0]             arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);

`protected
TK2&]AI^4@)@eLO<g4e59>G9X#P^39=c0Y6VW]\e<V89ce,=7886+)a3KC-1eOAO
#A2YH3I4JD0TfFZd=I.9DZ]C=G/K5NEW7_.IR];/&RD0:a@4W]bA52AK(b)c^@H2
=?Z>NR9Rc20=MIg2D#Q78gFU_4FfF]BZG42W>L\_?Z4TPR7K+\T(N93d+KNC@6)2
0-W7V44>@]9#6+-BFYVF4=gTQT5B@-QQZ7cVD]^HPYa,S7^=17_LW?[a]F6QN<U@
fJ=KcTIOT_GK?.[_1CN(BWQQ@QTYF^GNFXMG#Dc=5AQ2LB:+?4c)7,39,=6K)f\6
/-X1N:37MX8AVNYW]V-25<:P;eDaW.Z.CGDY?NTQTc/DW_6]FKE-UGY,)CGTO;3#
2H<6>SAF,Ve1Z+PdSBR[6PeZDIC((O;JeXT_XbIg1dWFM90>@=@LL3ESHGd0CBQa
0=+=+7R3A?X]0S_B;PJ7fBKC-?.Z&&PS-S0\<U[I8gO)6eUeE.^Z=&d=2.(A0A9X
\:P[&M=9<KPf7EJPKU@/L)c5,GfUH-5&MaCC?fG8FJ)-87Q]PS&HA<X0cbF)]Y/I
ZfbV,UBD0T.#P4X<_ME9?8NHLaP51f^(FUUCN/70@JXFaR3/XCCUTX]1]@K@Yg\K
([EE1)bF;Bc^^K4TDU6e9>>ePLGcea0?>=IA2e8g#W(VD884Ie1XEN(,g=X[).X>
a/OE(3#-c;4Kc7O-V^KXKVK\=4:McVDUUfP/HGYNGDg?6g8O;X4]IdY_>Xd]1Z;-
)0N0^FK#RGA[D&;g[&-K6(N1/^CA#a@Tb2P0,^)K8?OaGQBP6K,aFO;:.bdUVK<M
7O#/I3KRTb3,M+:43?S<UO;Y.]b:]B/+VTeV698)J,>J0E+I;?U@Qe-@BDF0<IZB
aR)A)Y\&6)+=_dZ31GTCAT3<(1I(4:Rb4(X>EB4]B3A]6/=?ZBWQ]PA]N+JJ0+(a
d;AeWE)C[]5F+[PGIecc7D8P3CBSEN:A&\3fd+0T(#9fHHXH/I?Z8]E6&K?Z;83:
)c5TN@=e&3S,C_W=+<77G40Y@]_&d.&Oa,XT_P,24T,fWOP;72gS;?N4cMNB)][U
KOM/&WA#R[LJdNV.)Q-Sf)YKNBBd7Z<gTQ@g.L?3TJ1]JACX-(6+Q02:3/:_ZMeK
EV#?>YGE]-&N]G^DR9Ra:[Y.NV@2b&PUA/OL>S:V?B_L:UEg]:VYK1P<X[<2fT?:
.1;,C,A+\HJJ,O)N:W8eeD#E^UTHJ_K7SI=Z[f,aFMR4?cF@Q]IgA(DCPQZEDL[&
^>XW7P\&<+V@GU<3WW3.J>VT)^gc/2.]QEC7X,Xg7g8()1ZCG@;>J]QI<G)G)-5W
Se2UH<M)(J[63]46e4[+_<GP<0]53),.#fIBHTZg/c<PPdNfUT[<CG.&GPZ@KK_a
50:V6#f#SET^XQX(R&.I6RcQ.MERga:1SEaR&N1L^3UgcZC(b?CD0/a\gKB@eL(,
M#0V5)2f-X_,\-2JAVdATL03Tcd;2912O1CB:cEdYBQW9K8HLF;g;4?]C8ORUVN\
dQ]aEe@C;M5W=F.SX_H3>KCK[L48@]X6E32Y1W-UABfQa?-M=LNf5G<FKR]C-bY.
0NDWW@75>V10R7>(;2QBEC7D,+=/UL2(e1N#OfaB^.J4WJcOJ<\]A>e8(?SW=9#X
WL?^C(D-^0TM=:eD@FC-M0fM5@+X9J&A4F;KVX)=FYCX8,g8a^C#KEa?E-f+7:NQ
2.7<JB&g61T<JWb#;JQLTP_<@VUX,-4gMb@(bPIJ3KE[;M0::3#1,0<01BaV=[^E
0>f+#/LO3SN<NQ#NS46^dK.gCD(;US@(LRdEabSg?@LRfY_2+d[HGD2&Ff0XAO(A
NXad,IJJ19\G0QaQd;@@BScP>O<RD+[&EPdTM-1PC<[Qg.H&e,Hf@ATY,@5JU/,?
8PbL]aG#XUE#S0J:;F1IN@:-[X1O<MP=:OABM247]A72=RRW,8><<^,(:^HZ3DT]
43b^_-@<4W/@OTZ\356RY7K>g+HAMQZPYC?G_CI;YgQb+?40(X9L=Z^e#>4<(2O7
>,8.1b\=^Yb?bAVf)DP^ZI6Ce1E1#4B?;c:>]@[:0LDdeMfIePbDC^_Y;QEeaaUW
[U@ee>e\WGRC&MUSST?A1&YaEBM0IWYETNAP/b_U<GVc1]0g:G#PIKe_>V34AETT
SZ8U;FVZeHWAgXS_7(X]<PWNQ^D_f6>+N8@62#[[TZ901T5g8.3)a(TY-;,HEL(>
F?bfRf+0N8R5]bEYG0g.=,a:Z6HK_GX70=:22D#aV1c^Ig@b#TJfPf4;7A\BD?WC
KWZ]N1<G)cZN/I5_#,,4a8Id#@AFb5(L[(JNFfY=]N-=7g+?>8M;<H>J[L_K\J77
7U:ce;eF]0eYcX5WBHcV7MU;8@dSO@C#^JcK&C/<3))a\g\J^;4-+?[^KcJRM94.
eJZE6X.:&7B-X1TR\Z&O&@88;_JZV_>DY4:ELW_==4A(6=\&9(beR)ED:+d-eGW@
#[C;MAPRYcWPJ</.b^EV4I]e0]G4U_-E,<-;J\[N>I;GGX9;83,S75L(+4_;<OOI
+D7O26FS1.ILM>0BL?+c02(<VUWe.#<H@9,G5Ra]T7]J:9CTXI.GBP;BV+Cb\_c#
/I++H6(2E)B5UW.O?<HPT2L20@60Z\(e&GXc)=<<_c[0@IE:5@.A+<N.JbNW,0Sc
S#V_I6VVYePHOJ_R(Z84LVeB(/>W,TE/5EgU=]KHXDY]HLI5ENXa^_<_2_@_3RJQ
7;4Lec-IQ,S4,-S[9(WW4\_K]gc_DGNa;#a1(HU^b-(UE,fZ=ceXd]@DGN<^M-+Q
SBQ&[EYX#^g5a.<RJb.c80b#5VdJ8/8#-NY=ET>K<B@)W&X)ACaQ^9,]-;ZcRM,d
B[_]C2a00A9(I^KbfLR\)S-H<d\c7VJ60I<N12,=8OVDG/K70-X1_?CMY_R?TY>.
bGGJ8+P\C&=R#MSg&2Yg>@.>.AY6U78#0WE/,-&-XF./<V\,^aSF^<PXD+D0[8N/
,#5VXd7@_2,d#S_^Z6QPB3IWT5==7FV;#f?<NX6;L05G-#L]LK6g+aJ[4>&e6:Dg
#TI:ALGT#IZ,4@@W_X/>]N<6(@c[W^SbKE]c@)ZXZX8NcS\b/M]080??.8&O\fSG
54L<R?-RYd4gKP^UbTI-9?Q[g1gOS_d4RMIWC,I@)F^_5YM8[R#,@Gb)P]O8>;37
OF[MYD=;g;9+Q;9c[XG0RdK+Q4I=_#dW];dN,3a649+902<5bSB5e:Q;9U&3(NfP
dI4M8&#)>+]<8Qg[O,@LRF6L-URdT<E8@)68O16QUa_Na&I@ELD)RJDd=>J[I1Kg
6R&#2#GVX&&4f5-DNdUAGF54?d<T9VSU^e@(]=I62RMPQ]D-R)DL#MRWc+;N5aHS
LT]LT?@(LB;c+H)6>1F&KLN12.KUZCJ&RYGUe^^ZTFO968Q&#3,+#K]SFTY6:bP7
[^::dW5_FF^5f(4?03D#XZ-gBL;QH0];[J@N=?M)=),N4OVW\]@##O]LO>V^J5cc
/C3X)M(.FgM5-M2((_L;UM1#;KT<>Y<_S/S)XW<^04LK:7UE]-cg@.?7=P3>b1U=
<_LLgCVQZ=MS<^5>>fR\LSWV#<C@O;3cKWVH,QWO<-27&_O9JC:R/M0<G[He04JK
.,4HP0C@4I2O,#<]Pbg1VLA&K;2#A0(AR)Y-_b-87Yc#BR.KFUA(E-;\cBP=PEd1
Y:J5c?<6HdF93=GDT&A\(01KQM704)M0W.dY[:?c=F<I=]D,BPD)8;41O9=[7H5a
O9PdF\]80S#Z=J,Sd5e.]dU+DR&P>)>U7CLe_V&B4D:GB#e4[JZbAJT:T,,,f\X8
e0H3(bATX94_B5J7Y7FPbO(-SIF3PMV(C&0&D?0)MBFIJ\OKZ[/XWI?1Z2c(BVTA
YRW8A;2_Hb9:C@Q9,</71\S.g&]+P6F6QTd[U1KNENB-63aDNRa]cU0S^^:O6B\R
f[DGNOc]ag<3c?,WSVBY1a2b0M>R=@3F6+4=e[1,8<PN7_R5?gRag?:]QW978-IB
:W[-/R]G9_U,+SH4\ZMDd#gg:/C929H(_TOK7e4WR02C?I;g(]#VKD6a6K:9IXM4
3.BP#;)(+U,Y#Je.[<c(S6OJ(V6]/cK^XRPR]CO#?G@gEV9>_ZC5O98W+P/FLV2e
Z4499X\Z^A#EO:Zb)PMbU9POY_W,_&(T6Q]3a8e85PEW\>6#ZQ[g@>V_^M0b;#OS
cH,ISX.A@9^D-N9b+)>TM<>LEAUE9U0UN]a-Sd4D?^J;@IACb-[76aP5P^AHF;LQ
U)[-IW/CLT,_VfLFDCJ[:3-5c^-(;^9@,4_g_E0a4SNR9e)9>U^PV@a6^dD#M1A.
c1UJJ2:4GX,?Y&231H7)&RXg_+ZAJ4509c\WDQG2E1-f^C]CSgP[\B:&+S7W&/HR
M>\D@&fG/5L0NU@C^=-:\O1@WgUZT;8HD2_71fef>8\>Lb1T>OI8g8ZS2B]RCCG@
eE<BbMFVKb0\AaVL/e[024Y9dOP,_#eH.7_&-Za;ICEJ7ZC?#CW[aXEM?1R[NP[:
WeUP)SP@NOa>U67C_<\Xg7b_RT(1KW5JN.8[]TS,)O6WZV&D;3(V#26dYD/f^CX-
O8_JFN>5dO&3.?DNB/PI^-+06M16-<QIOP0OPBN,^SYC4@Xaf?d\CVR>45fUWC]K
CLf:;RT-LM6-0I,W3+(bRB28C^WI3c^HQ08HcN+CHbFI6U9OZ]_DWQ:M5,aUYcD7
:7<6]@Y@1<2AaDRC;Mc)^a()B(<H7L-O@b4OMf,aN.bH<^[W(#O1eO8L?SSbU.UK
F5YD?6BU>F\Aa)Qe.)P]#XW<CRO9HE340dVAR.9ZI/]D9P;NMQTXS0CPF__VN3\3
=e3ecR1\:K3>4WfKKH&-L6W_WWR1K[Q[A^g=-Y)4HM4f(2@;acH-H3WeE,ZK&X^;
G0G7B:dN8SQ[CRVXTH24_[N=W.^#^GJ+V;H^T;.f+Z@64g0YF(-BdT(K8&cE\&56
CHcA/75.UBFZTN7WVCRS-ET#+NJYE6;\+aA1-/737ZR(8cQ4U+@E>R=)-/>OT5:7
__f53D7BC<883]U#:8RB8fe(TPDGWD&9)@(QX]Q<DNbR<eT?>&VO.W[A;TWYR\IM
c#PK6(gBe_[.W.\CWGE_+F4bOPHO&4g+D\4XCY.C--ZJHL\O.EZ0\RG#8E;7;<dY
.XQ2UKbM^N\B4\T#:)@Qd\=b?X<,(<>>15W@->ISD(Fb.4EXMY=.Z-Z0Zcf&+Yd1
F()D>0-;C)TDUIY)3B?+dB88U&(<6&KYb5\=@a#NE@0ZFD<+:;M]e;O[3(61K)PN
,[<dH\FJEMTFGfg31R0)B</KYMY2]T]+CA5?,U?gCVS(KBEUJ3<5d<O:B-(>S0];
^T[EB:4a2T#AXH,=.,0[-E#]H_6Y^[2NV890W)M8ee4#Xa\@>QQXfN=eK-+E,\AE
>DSAAFb<UWTBZ;Ef[0M6^DKI)8M,C6+Q^XUbZAc14[b@+)=],ULQ5C.gLT+901@X
7LWcYB_[(0JCbWd6EZ3Pa-eB96aIaA9Y.g+=WZEAU4\Q<,\E5+Q\NV);&+&a2a:e
/L\LKMbV2J#CU>5ZW8W.]DSL6YV+E4CU\=T7Q.T)=M?8c2C^T0LK2#S84g+;&A&U
gA#;(8e.^3EB03UN.KO\-B0AN\O[8e7b&,/.5G;T6e&aXDY2U9d<IG\@+V<.:ZC^
>AY+BSVe#U2&5SGf/1;B#e?I2bSGN3@8WbA@-ZG<AH>[Ha[.g7+f=.^QB.V>D7]9
);@NcYYP)-IK1ZP0H@fd=.\A-fD>YTNBe7Gd;4/]_.EVe(.WQE+30(0KVK.5\5dO
+Y^VF(0SfD=TfK1NF>@]00^d/8_E)WfL>96DY+@>S3e&86XHPf>9eSYXA@,_#Gf+
fLGX1H=C8TLQCbEICSd>U+E\/L;YGZYH2M;[_P)>H.Q9.]E2Jg2KV&]K[A-gPDgV
XaE@B[JN4c&,O\)(gCVUQg5<g^_&;cBSY^BXUCc0<[WBQR-W.f28#N,eK3deMD)@
I-21,3d+bNY7PAA:;&3NSO=H-G=Y08V65)1I6Z)Va?<4Z_+FdJ63eKeG02S7<HF@
839)PE?L5?12bAM>XB)aX_I#,F@IRL[IPV8#d^bK7U/_@IVAMZ3=Abg=WL681fE;
01G3BR\<6Ob:+)UGQ-;@@c8LBGf;5Ne-:VP:E?-\7@[)BTSW.WJ#,OH038[bBX-&
VdGREZFKWf>.L@8_0DBNbTH7;S3K#@,-C8>9;Ya.W(8A#MeE)QbdI<HFI0N2,-+G
-MX?XWZ.],JgD-<9(P908GD__.+76)RACWKDD7c<[GVTK2+)9UW-J[WHC<1:/P?3
9A\L7>2XV)Q#>0F26D#3D;>S2)E\85\)cb@8\1Y?Z[Y<1JXEYa>E+b\1HCFb>eH&
d#Q.@8/].]Z]470EQcU,0,WL;QZPA?]-KYPGDDc9e0A?NAOgG.,cR8\R.E@G?D^N
R4YUK2@C;:&=H2.X=c9DQ)T#C#?DVE34b,+fUB5H4IF7b@)UQ.D/g20,@Y7RP;0\
&#Q92D65cEQ54,+-(GU2OI_Q-LO4SY9@41@8P(2_e^Z8:J>@e=P)\3K90&24G[R8
6f7e;>d4)BbP/]/(PE7Z@bW+F,+Db1Pe@@0(abK1>3_](Z+.dG[LQ9aXB(f],?-E
7DaFR&GB\;MMC-&8A?34UNTO5GLF11\^cR))H_S,MZUXB#[^<N9&9+>eV>_EL^2X
X3W4SU1@_U5O2JXg_UMWX5CXPX,0C[\J3aNXQCW..Q7JK^.?Y<.+E]7Y_6K]/V1-
Y;8V_X^^(H]P_G<-9;&,aeX/TBa#GT,YB56BBNSQ-I7[\&3IVD@9LTfY\Da(PZO9
KPZ08MHC#<e,7+_;H:c:@N#N3;/NGQ-f))NFAH,6C(c?E)1S_A.K&e<VKQ5;S.c[
-BN+?]NR:T;A,Z&8GI=^ef,S_:?eHNE/[EdAQ@3EQ0:NW&U-5CR(2.G/8(&1P@L/
[-O0\ZPBO[-P8IC<(\UBd6Fbd(EFeNBE@MfTBgO3cB]@VBFd(fd8/=+&YWLIGab?
]_e9(?MLEga8W,b:ID945?\BV_6HY&:&:g#TgU0dPRH,RMRg+0+VOZ[;8Kf7CT[2
8+g8Xc9Z5=3cRK/eTTf_(;?+^Z&O2(/D]O),,1aT9T;(#PAb0+cf8T1T.-G@U/JD
(^G,dHE;H4-<6f<18-;aO>,)E06C[EIN.O/4O+/<R8DbW8^8DJ<^XJFDa-I#YaU,
U#K7WIB@.dQ[^(0)VV2G56NMLA79V;SKG+LIE,W:_5@,QgWRaC9#gL219(1)S-^D
f@R3,GIU0O#7NVNWJP&>O?,@VQ@3:WE-OVV\[QROe;,P1Q=HaO)>3LDbQJAEG7;f
W&+,_</_&]LHg+QR0Z>K#L#XQ0N\8;C^#PR/>#0)4-X:\ZCL7GD3(5K=L-2O2^NI
?S>/eXaLOS0RP/42EC7P]6/XCWW_PBLcF68;6J8E>6AMPbFc;CDT_82]ga_HN4?6
M-S(N>E;]+[HHMHBLa3-9<6,f;];2TK@Z:[GX>6U[WKZ#Ta/ASWT8?4JL)H?ad[C
MD3HQgYYK-53/?@:@=_:?@:=T.H]Pg2PBK4U<bIZg_XbR.>+9A\0,48?6VRK[Q?a
35?>+a=K(OY=d#f8NT;.R0QCLT776&8d<UN^2<\CZWAIe;WfOU4M_U-2=0^#&,/V
d7L+ZW&=/fJH;R\M<:(XFKN@<bd,HQFFTdT+]Va(-JUXGS5EKOV/NK)Z>_8:?+DV
gK]fg[M<^4d2X[U]7UO(TD(]/M+be9E>Aa[7Q9;ZWI1S4KGFdI@O)5G3(J)LW?MT
bPF<2BS7B>E)FIEg,]QMP?MXYTFFd6G=9P0#1RA?=097USDN_Q&YYWBDCX.XF:g3
H,2fZ;X=BQBH@0eAZ,G2<@D@a4D)I-FFTX,VP:9UE85<aHe21P2UT<;@_<K\+(Y4
)bYA2I@Zb49&b^A?VU\g?S52f3WA:547;MTS8I34C\GJ4,]IKV/?QMY>Xd&#3Z/\
SE<+>>^Vb<UUI]d)MM@F/83:5ATB/:\]ZZ4S^_dQ0[]/f3e@DK9RS&bX/]V#1;WJ
F)AN^(S&d7b<+XFN/UJLL;FV(df9/^_;)IVdAZHDa^6Z>Oa(E7(70C@:YdT^673H
@+K,?Y:gdTJOf6-U]U:)?bN^\/H(>?_HZRJ]ZSDVJ<QaFc[@9gEg][D+3>WA=2/g
-M3(VKP;>F5XY5@Z2MZ(^=1S8]ZWD=KP8>8OFd=\[gdR(fMYV1f.,K\^9)[D-VH.
AR7R),84)g.d\aYJ5JV6;,[RZZG\dW.f1F0@-&Sb(JdBNZOO5<2&eTT>FA<J)e_F
e3,>Q=O_/Ra:c;_-,]I&:H:.BY#MSd<-\&P3F&0SV>cKL3J?XE]\]BW8+?e6/-.K
@4CVJ?TIMd]b9VK0Yb.E3\S<Ie+(2f<a[GGE-DP/+)_CS8,6(QH7T1&T5MV\-,2@
4Y0=-P?&45JD2D11;5^^.71S5DA;Wc:eODb&1aK:=5A;YM,I?fFgEQ\Yf#Y2XAZ#
\9KO#cL#eX(^/&EP.),II;cVJ&Ka<+JCaZZ3P.cJ\J+@Y409RE,^FeU49)X8fdM#
;C.KSBBG;8Ief[+3V)2;<<@-8;agDFY6^_bXW(^C&?GebPd=Y@Sc=YLZgYHHRFYE
F_>14#CQ6,D#Q-X8^?@RA0AJRfPKJJ+]<YDZW53J(\gYadJJ>BC)+Ud=ZX>Z51KU
Jd][T5--f[^RWL78XW4OF4dd()N>@L&,[XC@d8cdA,<L8RMI?\ID(F-f&\4bZ1,R
89L^-Mc049DLRTWAVBR6#c7X1f\Q5dB&eg<aLUgHW>7I0-=]G.-5W[BX<f;#:ZK,
(K>S=eK104]^\(BBG_TXCRTZL14M.M#;;H2:@EE\#;4^BTLdOF.ZJ=11W4?VY_5:
2QJ[KLXZ7@M/fIBCA^:X2<GMPATd.?bL-SB.C--)E@KRGA4@N4;?,\5GZ9.4d::1
AR7XSI(Ne:#[WM5@I,f7W/La5J7Ld,S+70eWII^#=6=GKTT1)KOVE#bIW7Y+(g.L
6)7<ZPH\Z&4BNF/31C2FKTGRDNQP6T6E<;8d?KA4@R?)1?-@^)1.?bR5CTc@5\P&
a)ZU\OS+Wf5d-J.\dbJOHg;3NY2b&X&RQ7IH4.a-BK-X;5T6KN1Sb2C#WW7X4HBY
36bOfc2&_8LKY6D=0EJ=__2HV)g:2E9N96.UC[?SA:g(0^3D;5TC^-ECFJBEJAGO
.e5TVAOf_XD=[[XVXY.bTYcJ6WA]BR^4?5@7_eI;G@M:)J3?N_@W,d[8&0/Q0Q22
g6A;2DL:^7OD8L,\+51\EAa_+].EM1K[KOQ3fOGb@&?&J(\X=EXLDf9-IdT4^FAJ
L@8K9.&/USYU@\QUeCb_5T<DD2]6J:M\Q__C[JZR5(SIO+BgFE8[(]@4DbZG@-I=
JH.8M9.BaINT&?Xd2H-ISa+P7d4WB/N#O4JDO\O@1-0=XDRHQI7CRO@=&OB<g0Y_
I)@)GX62dMK5N=PeSCBfE#5QOLLQF>PRdBd\AdH-A</<<@HRYN86A\UWASLcA(X3
V]1\/6LYH++Y041</6f+dMN=(S?fBSagEN]S6K)JHVZMB&6>,\&PI/E<[4F-W]aC
4-b3K6)Sc1>TBa(I0@@G=;VCIKO89E\)CR8]f4FT?M9=MA^INROE+_\DT.4Af6HG
BTB^Lf:LQU=820M?R,AQRQF@c^ICYB+TSY,=2Z99ENL+RYAE3)>Cf&8G4cHf<>2G
<LQ[&M70F0d[7M]7\P__e(ST(UKK:2@YT9-fa@ZbX]UOG33;@TaD]&L<4bdUW,c3
:).e#1C?B5[-c2@#1;JKYIX:I8R)OP&0CV(FcTZG?JTU)B.I&dH3+0FV_XGf&<L@
Y\I/D)BfIEG+O&=\2^ZXeHE?Z^L2NMe]#\.?XcJ<HKZ[00@;CNH2LL[#5WR3O7c=
6FQ59+@VG2gOJ2\;W/46<c\W+TCgbH6FUSb+cV:)=1M>RN5,[8N?]U.QL+FZR,VV
>JOFY0e012^-W+[Qe)L\>C3.CWaFB^T.B<W<;P;EVCVf(I6.FM;geQ?</(E)R<<Z
CM<bcV4J#49F+ORgSHRVeN&1Be)+[ec,cILE=Y8]7]:c7SR8XW>cP^BMW7^Z)/>4
RL_IRgY]@0DJT_A<7)NCGRB4,[[5QO_SJ4>fAaOd2fc7dfFVY4]P_U]LQgKN<XGV
=&GdI<bATe&MGeZg^R.+_QG\O]O-fZg>>COd//c0PH#IB@])B00^g@g.Y@A_:\>;
GAHe?0G;ZTXM)C--H?P:TV)24[R6\TD<+]W.aWc8OVV;R]1^0d=/E++<QK<[;J#V
#cbLK2V_,5/2#d-<e2G<H:ZCJNB.T?aZ_?,e+aO/962(\L?K9cJa>@[7//=+@dKc
4WUe98Z-)9MdRY5JPH:-OeVJ=(?,IG1&2PJTSP0/?.>_X<N1^:fPY4gTQc:U[.W^
=fRa@7WDEK<RcZ.C]dObY@e[O0CATUd7:2]7c6^\^fT>NfB_W^QI00T2eY\-D&bH
YY]0bX:#\@H)RYBP[f/9/7?1GPfH:574NPOO#WN0:2<J#>dY\</;86-L&g:N9c<7
+#7E7D>D-[OCB<<)UcA^K;/@UQ86JL10b(:GPUV-YcceQ1F[3WF@R>LLbP<ZP?@+
ON)f2]a0gY>BN5a^1L\.0B=<0Ba[3X>e-#=>MfRKZ.86f#;.GgFT9^>;,HB,Q.>A
>N_\3QZ])9Jd.W8W2+?>6#fW@DCbGe-)g_@]2BUKQ3R@d-)F0ge4</>&&5(DUSFZ
-Q\,ZcL\I;P,ER4O]beUee]XFB\(gcOM>7H_&@9+F&WKOS]8<Q,_PNJ8aRe;<I;W
[5IUZYV?S\+J>M-5A?I&WF9O9a7Z)Z&TA=g7?0g[&-P-L(SBaDKEP]I2)?@HSR[L
#HaeDO+6K#39M]&Q>/XN^(J/K.)0MT3?A0QJQ_X5,AP(G:##2SLWJHU[6Q/3DD&+
L7Q?T+OZ-?4T23.FbA8U&0;RcdLAPQ_0ZR?RR-]cQP++Vd5<g1SU2]])?gC9aS^G
;dZ8c,&@[aEPb?X2Cf^#2W>eU/]NY)U5Z]6N(5/Y7;;eLPKYZ]/C5eK?(-9[RW-R
E(dXSU]EV4Md0BQ>&Y@b^<W[H9H)5TS].&PBE;d.If-(X&=#;\6.#8?\)/M8#=6T
e)PRQVR3\840\7C>/K-3<6,F\N1>6dXS3[DRBA#f6N]KOKT<0B6OB^9I\NT3WP[\
6=@?OOB;]8+O>WEU;2E=Y[M:FJ=)B<)dgT\f4(CWAD@+bXgOK[g:K2SX_UK>^f5g
EIE(RLJJc4;9I)_Hb>IZG.1KXfZ(dQa;Q1<22F)MMM3K/;c^WCSSU,R&=YTP9a-X
Zc1@eU&;<PGV^^^L)9=(aI^4Q@/?05M0Z14Ne.5,4+K#_=0cB0MeQ&bO9^>4ZW,a
HG.Jba-aY94IN+ecXJ8Q]]N\NP>>4cY6DH06W\L.c<&=UIe<,eX7c5YfO[aCK]Q0
(Y>[[QGVc;[)VA=dF[_e[Tdd[@)DeC8;bdX&\+[9+K7(VNc8(3H@/3cU(KV2X5dX
:W.54[2:Fa7XEa4<VN/dP3HbL1GMH>C;-C<XUdYVEN)UYSL\?e[Y>gV=(AE2JKJb
1EX,C-XIce45K+cLHAO0BaT;I[5NN_5d;@e9gd9a?YMRE,5bCV#[eT&;a^d:d0Y(
/3U]dB/?Q[S/g#XAJ-94/GNMcc-f87b&9GI]<Yg_aC65I^J8a/Zd:W,75)31R,[0
7.Z?BKU]BW+Z:>Dd84MC\YLMTLKX)ZF,?YO,@UOOI8_c.AC/32L_MB/:O(OD>=E+
<f_NC3?ISY(&VfW+Y1<0IPZGFI\YFHJYBP2c8V,P>\2eQ<-SH&_dD6MY:Id/2U#>
,(cNTOZ_AZ+ZP=f;I8c>_8APH<]9NH>>L:(94f(f,=JSVK]3=UK.L/+.RWJ5[+\]
6ML)[1(e3b]N,2<M:QF;UbcTf6Z;Rc6:4C5U(,4M=L8,KK^2C@=KgHg)2DDCC4#8
4RQ4;UFB@C3DEg\&9N=Fe_.[=-b7]K^76RU+L1N?OEXF)\W9_0d[fccIB1J=ILD9
fL+V_<eYE[ZWc8R(U,M2SOfT3TJV);HT7TY;;C?IU?f]A/:@F\XUT[g8]AAe9,^Q
>5aR]7Z]eY2eNKU2-ZH3df#]6f/DSY=fHI#7HDf8&#^(K22aD/UbCA0gM8XNfMIA
BQ_QTWTM)VI<Fba0W4.O)a,S9TV(QN>HO0MX23X^&93FcZ8KT,CSf&(]3QHSQfa)
c6Q9A/Xa2A6^@79LJP,8U0De0eEA9_bW=9L1Z3U\4b-aPAIM1U7D55dQ]c7T(b(R
7FUKb.APeGI86X;aAU-PZJD,dRd]<MPX-3E+d#NOTb+cQ+-#\..B4b=G\>dLaZ^/
3I[aY9bf6&K42N8GbRB9;dBQUV+V)1WL6=AOd:Q1d=d+=/GKSS-6&DZdQd^V^J7U
A495NSMgfO>Q=ZLU.L3AFF@eW#)G8.,0XY.b\^BHaR:Q(D6aRN_ZYJ)PSS:]?KKY
OJDdE,,DEM^dcGC7caCBbZMf[GgJ9-906OR-/43+;XKNQ1OdZ>b^A>3,9X^-V)a.
F^WK\<18a##5b&>F^2JO-;M[Z90UZV[-@TUgY94Aeb=O<EeYW-b@OI=]S0a3W<fV
c#Gb3@PLNbP:8<9JQ9K<J0/+@bae@<aC,OVZcXZfd5<5>_.(.eH:.I1M?XBI7M/>
)SXA,T^>FC)SNYMYKO6OX=3UZ72cF4]C=<DY)e2=\7XX_8_3EU<3,,/a8>R;ACTW
d2&RU;DR;?&bJ7Qa)&,BCcEQ=4L54X?TQ=&=6W5)N3J/7/A9=MfLBO[Fg)YR<@=?
UO^J9MH4.VFf+;VV_S3RK1EbDcX=6\PDf8D)CJ8/+<0/M2,S,1QO-be(B)&\M]aZ
);3M&YLb.)(Q-UPD@-5-BT#&e.4<AY,S<c_4Wce:(3TUEKcO03N2H)8IWZ-#?+2Z
<EY8Yd1X\T\R6)7UX>K.1&)cY,E[AJe@_B&);c0]^:Pc?2e8IYbX^;\KePa&E883
,dNU\F6=&?(T<FbM0Q)E@^)@Ge,cN[bfd(;6+6[V^(R??C>I.1#)[Xe=DN,g^Ea^
?406g>:f,eJOCGPI#BX5+);.ELI^6QH36BSd5OF0WQQJ7)W.C>4ER3@d#8K&D6EK
K(9b#<6c8U)W^\)\(2(X?1BSDL:,LKc/5\QR91E=[>XZASKAgg[JPbTB8I?J45OZ
[;J+F>VH_+[@O/)<Rb1g,WM<P\863PTUEdUeK]GW_cWc^QU061\3&O.N6(8YO<_8
D(VG=+^&39.5U;)6BZJ9V.X4,XUNKZQ@7;dFQfHIKU47]^M+X]#ZGb\?18dV@HUT
CaPX2-gC<4B#([/ECDKcOFN]D45E^ERXcg62?LV+:M-2VT68(6NM-P2T^59e8.Ea
>J9:(@+L4Ie3gRW6NSG9HD5GgM-e6[6^A3CL^fXB,QW,V@I8-Z@a]_)G29d?_K<(
H#+U2E:.HOG4O7)a-bf,>VU78T6^5DIS+XMdK&[7U[fFGL&?g3&E_dd@>?,(b/YT
IMWVDA)\8=:/8FDVC[]NeNeDR;U;#7BM:?U_NNUQ6#Zc@fe,Y>)528a0<<]b^(]6
=_8)L-LCd5J;XBE0CJP&\1&55#=?6gJ:4?c6gTNYU(RJ)GZac942Q&1)0Kd7]7Nc
FY_Q(+0/2A?OYSX.8g-;TL>7/J>),K,7QDOe/fVZ-=ae:9,,=.HR4eea(Z?[_H&=
Xe^gJ..gHJ)=QWgJIAg_<XQgbAVK:g.PZ?YOa5H4B_XWdL.<GUgW<FALUN;C<)3W
B3R4g1^,a?-1IUXO=_<JX]\Jf(8eL6.ZEfYZeN2T024eWXd:M#PW;75N4GbJU7e:
@3L0OgME2[[HRg<<>e)_DH5.;09+E_KbVfO.L?DLH-X(_fAg6=N1HFS#DG6bM@aD
9[7^HD0;[NAaTQ[KU6=W4P?#]4/-A8A,:9.2J8R1a;48HKJ#AWY:5I.RTI>MMD7+
P7\?2;D+b(>=B^E)b54J>bX#^>GaHB1;,6SZO;c>(=>NU=N:\gP4B+-KIRE.8UOA
L/f(Ff0W&R5@V2F0@4gW5g9B,RZKY)>Z;I^#T<?GAW?d04#bW=LOE;Rd(U<4c^_,
4\7MIATPc0d,_dKcQP:)V^=?719/M#ICOEXe^gE9M(Le7D/Z\A#\+gFGc,929/#\
,b;]SFS)74YH4a?^AMa:dKNA<P6Y(K@)OUN8-d2S;;U445EJVQMT9<OdU5@,6T;T
S?/YRNM-P:bBOF8&_Rd-GWf6&AC,5/K3<_EF#T?VV#7a0,>cT:[1<BaO\030?&)R
dda6706=-(+NSf5P:>J+G^8@JXVZ)^D/EB:^E[M^B8(LF=9fAaEPLe(5C.K<KG#[
GVIF:^X[7B0+IUCTaDeUCH:3@+:d\O2Tf&b;-=)0B2.7d)IV[1WUV,^]WFS3X@/D
EX2,;&DMQeQAc,ZBg5/\GF,ZcKH4Z:O</0WdQ1CX)_3ZK?SULIg<#_SZA&4a8Zaa
0EY4=U(aF,.AXNc2E.<9KVe(]7QZU\0-W:6\XdNb3<gQH?+f9Sc;/5M75/)E21JB
FAB]-UVK,88#EXGaU=fXNZ:ZaFM^6C\4J,KfLCDf5A31JF@FKIJ<JQH.R=Zd6-;2
&Y_/Z/A.c_X;:9V7)MI+QV?9Xb_DRZdFTFH<bRaYK[U7;Lb7f<K&<e/_fJN>,[48
S>Cb.M+ZWAI+VUW2.-f^OIaZ[:YYE92PE[Q:RVc+)G2?Z=RJ?Y,FOfJU\+TF\e_(
>8\L)VO3IDKbHN)S\R#/E&IBEe5VbOFHc4.:<ZEF4P<(EES=90e:0eDAZ:f5gZ#F
LB\-(1)\<.7DZ+\VV=IP]@DaTZ;+]1F+W<X68;M@G43X^./W9=SXZ0XY2#E56NJ#
(8=^&\Qg+)DO0684;X.gb0EY[=21VLgL^<:CY2WYM/ORADBQW[-]Q#3NHa>6@T-T
PPYdcf8I1QfB>a9Z>3_&4KQ?+^Sb75D&g/aQ\S:V_QeaOXA)Q+(f^fS@-+gNE^WX
DAcP)\3B5OFO=V&;1013fI_e=c+NC6f=I_aXP5Xb(N5a]FIMV_6QaHIS8R85,A1]
NQ[JJbb=a>_0<X6d+1F]#ESPMS\.-^g,fV@FCbC<HR(#X8EXaT-.\?MdP8SFXAO/
BJ^]6H/O<P^UZ>D-,a@7a04B:]\WW>8cX/)^PF??/;PISY,Y-YG^f>S_HeU>/ReO
>[8[_:,V.B=M=>LU0G4/##^Iba8^>=KO6J1@^Q>-4PGaMb>1\O^)EF+dgg/PJT=R
E-D/UTb\<G5+D;79Z/?6daV#9DY:U\B60)dc^,PPdVG=G2+8+5g5b^O+CY7T_X#O
@1fR+V:.(=HcC)NY0gW=3)V95R]/_NZ.9TPg0Sda==B8BGV=g9)a>CAD8CB8c/-G
,9KT&3Q>MX4?TI-7(c\e__UWC;)b3YdTVU1\;B:2@CBQ^.L;bgG6H?^GabCYVMRe
g@T02<g9YIC=@4UTMeN)<COMC#WW?f@O^B>JW-\:@3A5[7XP,YC^ec=6W)XeG]fW
487EW;cJF06]\^IcLLf)9fX(K?0b:;@Q3]e<L9):eaS\c63&Q\?O63a1TC\BS<8b
ga2HVaKWLd:_4237RGSF8-6#E/:4e=R-Se3NBAE:M_V-6GK?C>T;LSG<9,O[Z1/R
fBT&dF@fGY5APdGU8]3;P(Z.JIN[Z4.Z(8@aVV=#<_VR#P81cDW72KQ4-NZ>9:#g
.XA(WYb]Z<G1//U61;JIB#2fO6K_6;:.BOE+/F<B[O1\VN9U&>L-YDO.SZ0aUH2S
#=/Y[e9JH)/>cR&QHB9VHZT>ZP?YNMMYUJ@B9C;RS=Bdb)K>._WCY.A0>a^)F^+f
+U&/--Z+\>P54#I+/?8/EYcgX:^VbRZ0RVUL[AI<?XDP]<De=[=6fUS[Nb9DgOI@
Q#aLW);.>f8QFHK\Lc-.P(4A)e;)TR2A@LeQF6dd-g[_G.H5Xe.UdAO+CGgB56@V
Z@8Qa.1e2IX\R7J@@.g3S\NI=,R:6MSX@?FW._DgBC9d1b4Z&_RPEJ.:LAXS4aS)
efG#>ag()cYSE^,3]EFD3b_fUXbg+/egbDNgWO.?@g7J:0UKF@X_Z^eaC8&JILJM
,ZT,LMZ[6bZL(I8Z=4\a+S=I77T\(:^.?KTC6aA\U>[)geJ>F53+[>XE?4:+4^?2
>3MJV4AXVcRKJN,gT^,MNc@eIRb)1^e=H-GVU9N-=;fc3-&fB:Z6=(c:faF=J.e/
ER(;]G?^[0JZV)ed_H1.gOf@&>a(425R]2=M(Z3QR>-)K]N=[D0SaT\6\]=2@J3:
/)_Gb)1]X:623^bD#HcA6eNWW0E]GWW/8bEK#8FSDcA4\3OaT@fFCHg9C.^R3C1[
OO5a/22D+,+LW\?f2a+3Z[9.2HTW724L,/X7?WP<PR1&9/K=<6?7>T1OSSNEH7/=
S2fC=2DRY:[WYI,QZ-LEe0g._QZN<-M7V46W^()VF^E;f<;QH?)>-PRVC5^L8U9E
GJD\_+M97FQM,Q\L@6b/ZGgd=1(-:F)8S_[OZb]2gXUPd2[2Pd;[Ba)CF0fTb)^-
^eYf(6@?Q4A>H=e.dN]f6fd[5GUIcBH67T)\-gESIN4?BA;3DWYF[Ba+F-;HFR_3
\f(3dJH]d99BB:PTEIO<UXdQ5M@@g@dQce9=2eN,P[CEdG+P?#?W\bcC&5_VIM@<
K_MW,ga06SP31E\QfE#8F,Y6R#+QTXc_HXM:KKb:;-,3JcK-5cDYTO(&E/8XdHO\
d#@O??=L=:MSg@(2>B^CHGG.g#b>59IaAHB^C/+Z7Wa_B4+^@5RCZ[?^S0G3FZ#a
5c,g1<#;WFaYHcG=20FFH.[Yg15@:^=\^=]E:MRg^H2ac)61:QWDZCe5&dL2>6=R
<Zg)O#IV_EP?(L6]K_L.,(N?ec#U)aC9Ba3P]/>RIS)0KP14S8P:4,?LMAM=S5(I
3[T:40[^,H_AQeIK]^XEc<\_#19+L98S>521_?dI_[9ERbT>LM?FEf1?28,G:dM1
F</M3Fafd:@(2abXR_@D0;Q1#ZHDNJ#YM\)#4CS6:MDG0Ff+Z\GXd]DZdG@3.R=9
cB,(,N+(c.ZafVVU?22M-EJTOb\Z?Z#;MR\]<P4A9(f/f_YU;1Ie0G^c-B9GeSeQ
_a5#T8&Ee)V<@1_+K3-FF3VM-@f?ZC=RR4?48X4b]L=LLe#>58cV??A;6=^(9(?T
8B5dAR7;5&)N:a=6g]9>8e.NH,dQU589)f7J\WI9+:FO/M.CK)9XMZF;8gLcV4Sd
c(KcWLRf[I0CSO3?O\(HGVX)J[64FV)gICB@ZFQ<NDKe64ZHdgZ>:#J13.:ZC^17
?+8FggK@,&eZUII,1.)HcTB8X/(fbb51\=/eKAe-8gONd(9U.>94C04b+C9,DBNZ
AWOXIe;<JeP49?YQ;,VWU\#f\5aEA4b[QYV&+;,5/EW#eU<JQHJFC3@3]Zd2O=EB
QWIEB+DPE]IE]DZ#VH816(TY;0Y/>4UR+C6a9>U.E(@?aWOc@&7#TVZ,)-)9U2\4
86;&;,>Ve>deS]d.0Ddc3_P7F5FNT+6DdRF?gA.S8ZF\Q9WTE8-SH+.,77Q&)=\a
FP?PF#M@8</0M/aYD]/2TWGT-X^?T(0Oc#;O7)N3)9SWCeP#d&5[SaYaGAULdKC9
/)c4_X=?LVN]0)N<L7W0?^HTKbG=5RfV(-]@5MNF<-31/e._e21RC[fIRK6WNE9E
>@/HUb3PSP@adPMR024>FR-89_LJ4NJ;f\&1>0MKJ#B8JZY0_HBQ]_[JG:#H_X_6
e3e)@V[=5(G/:D:@R)5U#32N^@:Z#+.E3;R34PQd80XJ\9NBF[3;4a5OE&eS9,7b
1F.Z3RDY_8Y.HJ&-R58<]K[d>?I<MR<#1N-TI])ES&9\-N,@A\5RUF_)U=3Hb[;[
a<?]Ma/CATF\&K4ERN3INHeQT\E4Jf_-1D<NA1:>/Pf@^8a?N^\c2RHSFKE1=G/+
LZW70O#FJP1)AA85?&-1-cGJ@_C-7<eQ.P[>eda)bfLHEWYb]NY:HZ&,&RJP_T(F
^@3@E#(1(4c>V&##7_L&UFX3,9:5)+G4F3L)0)H-]\EF0?6gB:L.e;:J;J4;P=8c
>2F)CY(&1+bD@G(fN7KX8&L/df/?C<4#P[57N]NLDHKMN_O:SWHOFc1)aUZMMV1K
Uf4,L:P9(SPDf5f@^bLG6eUMEaW;8/(BGC14(EcXE8T73P/ELCaRed+NP=#Z-@U6
/:+-0ALeCZY=MI-<V^R\2:(E;5<:KfcM@;4F,<74Y,XM/;6P<0ObRPW@PZFB5cWG
#0_T&@REC>XbL<fbZ9&OV99dfC4[^[Q[D#:T@b0GK(fc;S1ZAeW=U-83@XFMVd-M
M9aMO])8<Tg>WDc&_WZf=4W^#fff=0]WVHZ=23Ad;)UIY?H3dF(ZS?>MAQ(XFe5Z
_X6[I@Mb:LDB1+VI:(X-1TP+12GURc3NcKLgdYQRT(QK8AD9383T&],U7B.4G=H1
93&;]\3#a0<Lce>/DL0&B77WBNZMC#LgZLUJSdfQA5X7]TZVaccB\Qb5,<IMG;6R
e^ZgGfIN4XV1(dWgA:LF(>SF^N(=C1T:TS>X[Jccg&,YVG6AX@5UgdHDZ;\VOAA;
W#[-TZ9]B?P0abPEP#0L(acIXFa\B:60g3V6[(Ia:_b\J(&V\01<#;E.E:UL+U3W
3HJf)FU>)a?3]c60^Za/R2eW221&QF[S-S9QZTN)g&OVOHWN<;;>211^G--Qb?M9
V)FR\I2#_;@c<3NUeF64,55.LIJF2)N6T;2#Q/Z<PWVa5ZZH3Q?W(+U/;5X.B].=
Iba==+f1fScKSD\K^J/;^,FM1_]>IJHcgfg44PT<(dK),/.VVDR8^bU4)YaaC1A6
S]LY@\N3efL2eG>3CU>\^B-R7^aOeLe0[;:9I#(PCF:EHf?687/IIMRLM4NaTH3H
\XZ;3.]P5^B86UBKEfVHP^IfG3N1MXHf&gX/4K)K8<a>SO@e1,\eVaCMH6]H,L&Y
YZ?d#Nf0Uff9;).;gd@>2.U_Z+O7EZ1J[De^K:QN\-V2D0c1E(_FV;P:7NNANFA2
\0VZ>Y_a/.4>-[9RQ.HfKI66/6?B8.A>6aXP@<eGCL;=T3;TI0&3?F_,=b&>AJ\c
S54_O/N?;O-247gXUUU4eHc7)2g:[;T7X=4EQ4[F&5?^)V^P(I<O#0IJVJU:O2FF
GGINA1O>H3DP#UIJN9;FZJ069L#VL^BO8;9F#HM5Ee7YC5gX8/W\?BXGW6DVgZ4&
YEB++3MA55:HU0^<4X]1##@NAU=5P-CQ#C70EZ=UFM&bP7Ld]g<Q:WF>Y&F+9af1
(B(a<(9c/[d3E)&7a-fe5WBa29FgGU743VMdc^HETAM38#^)DMT9PD[QO+8MK(U+
?^,.(YTOK8cdZfNU7FLX-6M.R:<X1)[<W:J;A/QfB7f62&(1KceKeZ^]OIGUVOf8
EFL8O4F^#d6N&PbMP12CRNg2+E_e:fD]GY7_OQ423;6IX7C3AX-eN_:CQ,B<HC;3
EX&IV^&f+c+OG7L>N+C].J>@a-EL^.3339O;16&Z7OWEMQP0#-KS\g#fcbI.(^P_
3)+NVFDQ0[g3SNUR=1<E?WJKa-H+NC17:=0Q76L(c,2YMNAU(/aX?0?,W>Qe?,FL
K4dWC6+.H0GQ(aD6.;8OT:4IMVaWEBb]f049;TKfKG:US6:(WTAF21BG2&_>^\2=
),V(T?^=(,JH(A4-T=,9:OcANWb>;#IcMAO\Ud1C=K,5M&]&EgPZ3\1gXNU8(@bC
OKSOf+Fa=0fWA\+P6&7_f3f+2I4R3I(W];@=BTGHfNU6XI5@SS7f)/FBK5-ADUT5
Yb[65UI<O3-/G;b)49GZ6;#649c;C31)&FE^21L8VKW5;PJDV1VU4E9979I.AGb[
^4Z\:d2R5a,^4G+JHMN^QWbbd2??.^EB43S-QE;((2X[)#CG^69^F4bA&^11;A&7
aFR:]5N65K2PC],PS:FEF(4LBYgPR[QT5K@a^fBVA.;P?<.?M&7Nc]::P\ca^/BD
,KS]XH@@NKc+;OVPZ\;X-B>cd959IGCN?^b4=+6/aTbG7dG:(EY&G.@(H4eZW#_d
@;8(54RE</\@.L<:RQC9E<WOSX#B)aCMMgV5f5?Re)\T+Y<&9UfG0@ON3[6-+(MV
#[+D[NN_ULX8W52HW_[8(;OgYR[H0DI?cceOc=X(0/5e7aN/UEK62R74Y;7a.L][
6A;B\3@/<cd_X//<Z5&2?0;S6;Ee&_2^47.4JaBK&Q</3,;g[KYeFB9Og:JZc(Q9
@a>9@K^=bdAK-G9CX#@O;4@Gg#dZ)d+CU2f[2/NLKWQEL95Pb#P1Y1<a#0bIZ)F7
P\:O_;QOU[?RL,2Z1:B_JA[->e)c;W3=bBS:>,=DeRNc[.?00:QCN,YY5];?9(dF
&#+QC.PST2Z2eHSXGZ>8Z:[^6GO/(8C=J?S>153#/XQOENKYOId5F7:GGBf@+RH;
IXdB.SDD>+I8XDQ(ZG,B2Y3&g?,B8H&@@BW,UD(<8)JW8#F[Hf2Y.S/0d=N/3g=5
W+b<2??T92=TT?b[J9RZ\KQgVV90KfHWGa#?V/5?FeB+:f[W7<F0[8L9Q</BF2BT
+>#U8cYfRGX>8@K[_g>^SDW9;->Ag^-VN:0)H66:)Hb_ZT+FV]-;4^e4>X9Hg2ZY
79(MM;>A;PX4=N[[6bI8M.<<e3@[6cB5ZEYQ75d9;+96W0/g&)OLLKZ)f?(T-VTd
I_>fL1GGIF7;M59COL7H,LNGdf(N8./7)AARNJ9]eAW57C@6<.[?^PA57;V+_C_<
TZE]L)4JL:T0U70/C<M;8,=,7:(F-K[2>3&#\5[\5e_A]d_)3G8Y+4S)&\R:S\_6
2+3B?-YI5)3^2YMIG#EW;5]_b5;G.YB1?V4[2P@C=0JdAR+Ab=JH\G5:9:G)7_S9
9407<8F&-U+b,Sc^cV3SgbEH@3/>/?43@N3QBfY1T@4f\JDOH^N5./IMUG4GM]K\
VAMb&NgWA#FgWYYfEHT=(=#>.D5CF(OFP9=aB4#+?>EJR>X2;2@f+:IFZd3?<_@3
S(Q/[&:;a:EA8fZUAF],#b-IGZUf\bL.N9a_5B9SYU=IC;[^S&LFPX4&&<L_?C^<
M.E#KM1&QTA;7IgQd#-_Ba;+KCQSB4(>:\:ZQ&L/@Y9+9_2FVX_#[I9_/5SJ_GEc
#Q\NN=Ye;>FONPRX._9]:#(CLZEOabgN^&50F-1\ad7f>c9(1A.a2.^TC8957GYJ
=fPVP31#c83]:P6M(69F<eI?[/\[WcA&8L?,?=Y+F[57g0B3c5.0ePaV4OcKW8dc
I,8]<7)QQ8f^[>fO?a_5H=LHDY.4W?&#Vef@&7O]OQK&GggVV:O2^Ff]E#2HSceS
_a,W0&P6L<Z8PZ6FHTS=]VJ@BRdf,7S3HGBD..H5bH()4(]gZ_E8F#f4]=9E:B.V
PMDFVLXNZ]5)-#9P0AD304O/bdJ:O>d82NQ(+2a\4Ta3-fA98WZ4EN+e]c)0&;Fe
1R1<V\/ONdc?1#fAH87XR^(GPO24Y<eD=]?I=[Q_Q;[RZ)ee<PV?AV,3H((T;X@&
7V#C01_,EP8D>+9@9/a6.7=I,+C1Gf0F^N<MeV_c6J+H@4JDdbT=&O>H2_&I,RGS
bb(TJg=C\]?Yc3-QQAN^1-2)CMH+PMU59HT=N=.8Y/C7D_T/09PPR.]fQ(3I;]/I
MTb?#VXYLH#B-9[JWF?XULU>1@,(RC#P_R6f/:VCP4+:Q\6a)fRGBT&bIJ8:4>^Y
2Ufc_N--/d,-1c5ggQ^=JRODMea6:6?9@e-e#FYT46.3:N5e0.(VcS_O>X&^S4T2
#S6&KG988)WBfL)4;5FW76K?KZ0VD7A,XC>[+,G=1/5bXQFYG;2/3KUReb)g+a=4
N/\Q3daJ(VH&T?7C-TN2U8.KTMJAfOe3X6#)@<RN;V]LP6FVB5Y_^E6c?6>Fd#.?
:GK=Wa0X8bS8>U+/ZQYd#g>aI3==T77c9>JA8Z]e-O7EXf3>PNfIP\1XM^F1@,U_
:S@D+FW@0D:)\Q2.HDXcKL;621DR1S,QKM@H<6<(XZ6/Se9WHUD,,+>@T#CC07R:
Q,58aGJ_LH3+ZJeU9NBNPIAL8Z]]dG>8NG,bS</,Y+\_R_WGc2?AJH3O##L;QL&G
0:0R2R<;BdEDdAa9NR?a0]FUO?K2]WB=&7Ff)??MefAE1\711gfX-8bgN(<E_@7&
Nb.27>[a,_8F.GB_aA:GLJZB[YT?D2PMaY6^EFe11#?/H7GdbL:;2=IXP3L3#X(_
[e=bF-NS<3J:R+@UJTeRWYQ3V+gR-1(G1fO7L=>UMg6dg9MXdEUJ=bF8\/XP[1(E
M,S;ET0L<PZZ)>1Y,WF-@B.#g5;1G<I\a8._4:=gL?J7gQPV&28;IA.[1bW]Af(1
2,QPMJZ)^59Q43.QKdQ]e3C,^FgV\0-OD3X<36:=caR[@J8047&[Z&CN]8.UPe^O
daV5/b]P;H:NS;fC1O+^/;##=.[[F>?L6)J[K45\fJ:,SS0F-27Q_b#_>854>HB:
DTePd+7c\Dc8;]ADLQa65G5-66OX\K=aYZ@H.D:Q_2LL7Q&HDZVNXdBV69GL6QRe
Mg+5UYT]Ca&N.#Tg:0d:<,7=f0W5eM1?[./J59<=KHU2<_53C_^.COH#FBCS9dXZ
QddL-ZM83+T48W1\f[=IP_c8,eFfM8VB/65Z\HLQg]S^AJ3_5PZD>2U]Kb,gc&Y@
>PM[F5Ab:0Tc?b(WGe-JMR8d##-f^,L,9+RgcT-5]7B.>^LOF[/Ra-eUXVc(RaT8
&=(,[e^5C4RM(;XdS85+IE.DeN9C-39LOPHTFZZD-QO0[cW3cfcMY+XDZaOOP2,b
-_/W\.H-O&^V0c&Ie@K?2+ZNXWFQ58HNS/bQT#7G(\]Xa#T]D?-Z:VFN18ME.Q)T
]@<1eQ\4/\,7bQX[9G?)+YYZY<WE:D/ABHg74fGcd-8?68,3[KN5[DWH6[\)0L\-
.I4],L7:9B^MU1dMY-P>##5Y+EOMFTgA<OV&>.OQ&-&9b/+3eK@+2776HbD\Dd+S
D=&Y^9W]^D56=-S6PHT2]:4WQ,_,5a\NEa;/N.BK-a>Pe/,5V6S_O8[ORE_f^&Wc
dJ3E&+RZXCd@ILI+(IZL[b\Y]3ZR8d+4HE85V&Z_[_Q4AF<5B]2:),]UaMON&6#C
&LXM4/:U#S?a9LAT3(#J0UCaR75AH,NNH),D)]6b^VX<bd>I>aRCKRN)[ZX]JfPQ
,Ce?#6bDQbY/Y<_PJLd8K<bB:fQ/[Ke#-g:a86Y#PO\Z@#aHK)8f<f55d>?.)C?b
FbCHbfC/fI>\7Xg;9a&^^(YT\W982&0/FEQ\<K/c7S:7eg>^IFA:CJE0=D,DO1&8
>[,\K5DJF4FH^4^(LJ^F92]<=]R62a?._Me20LZGEVe##c#0F]M8,+VH(3B;FIPU
BOQICDNKD+Q<Ye;7D]Sdd5-:#4J/RZb<DO)ag^a@U=A2\cX,(G&e)G6fbQeXWHM[
NV(RG0==2;->)].Rc5A7:#7I)V6?<0e,afL&C&c)W<9,)B>G@e>f4#:3L,Ca_6]f
bD<.]&T7.8V3+A:\N4g/_ES+afSe.Z5;;$
`endprotected
endmodule