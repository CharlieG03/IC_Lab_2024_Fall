// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"
`define PATNUM 100
`define SEED 8721
`define CYCLE_TIME 9
`define DEBUG 0

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
c8RE2-^_7CS=AT]YFYR9?_^[b-A5>2;c)[55g4dBVeAg6aNP.)@a0))2_HZ[?YQQ
9cCZ,S0=PH/S1^\aWQ,5f7eg8,c0UVI&_g@GZe.3Xg>[SYKN,2(R5H0E=9Yb@L]<
I4XRY8D[KW0fTa8XDQfae>&2_IEKZ><-AO<A?7cAOF4L]MH(FF,4<=;QZQ8IWVKN
DH<[T4G2RK5b/0X-:\4N:bJA.=^O>cf_-DDg9?=UA+OeeR/#V^K)T?\ZTZ\X;J=/
(98FQ9TR580<#H<_4bI2:;a\a=-&_:]2O59]^a]=AULYb0YMHV,TZD^aN:fXG;O,
V],5\W5H,;Md-79UJf:faRJ#JU>PWgZ:=K=6d[_[X[g[I4,E@K<aA3G@-YgfDGYe
#>d#S.YH48+E<Tf74a(XDLYef59J9D3(;X3TBa\];]70;N#d;f;[M<cXD3YdXeg[
:WM+9W1M?K2LV0Ya]8O@.:(g:17/Q1#-O)FM4#?=G9aSQa/fc,88<5.L_@.8?M/A
5FKG<O)0V@f(b[&PN_H@d@BON\[aDW-W,Pc]E4&>c=S>M9OCN42fNgC8X,_#Nb/&
5TJ;2BF;4OO[Z]aZ+/G1G1dfMbJ+)Ff[BJHc;69F=/EMO7:A>PTQ[UFC7:Z<T1QJ
afK5[FX04>73SaUF(_VD[GI9>GE.gB9LFa;S.9U47<[^3&)<VHC[P7V/T^]<Z;>6
8L/S>/:5[-a/+#DF>:T]0_DW_1;R0_-ef1Oe#8KDOd/7:-/(&aP?G?_>,=f8;]SG
c(IJ@d-KC[2COeBBD@)QCW+]S9CZ=?Z<_-G9[WSB-7e\(UF==DWS^6S568aJ^adR
59B[_K0b4Q7,.GD#;L0<fRCFfbPY3/C?P+CXQP3FEJ0KJ61<KSb2@+TD+[eAJd-b
-V[WVgBTgI\:H_4WX25]PeX[[GI++-2J5K#?bIW=>?=8.-J=J,J#WA^O19^ga0(c
@Y)ENZ8FV=H\@VDBVV9+Z8Pe7;[fO2FS_G+>MVYS;_7Y[\#[G_8F3IH4VgIGAa<b
B&TAEP+BX67^c<]/^:g@;D7HP^gg1>QXKY8M+Q/MOPE&eB4-2GT53/A:C_JQ35]a
-a#-):WG03,W>P,[^Mf>/AW\X6(=V4DCE7VVI6aAfN:4@Y[b<b63U6V3JWVDP#S]
=Z>Fd2eMb535D.^a(fdCAQ9#RTgg\&JRKAA8W>T=#2CN_C.5O-Fc#]/-I1V>O<Ga
+=g4E=^/N@WWS]1\]:Q-.1EW#R&K]=@YLZXNO_\OF>_,F8ae&=VVD2:-OT>-I3L+
C43P4ec^e>9Jc0PYb^6N4KT^eM+1#8WSKCJEQd2EI;6MVV@_bSeZ2+DXaN7TYUc;
)?8AH,8;S9.;3U6G=DCE[I?:f#(W2F&:H9,KMe=C2XGKRBf1IVe25PDT?begS)8S
5-#Qg7QM\#H1RL.:O=C@8CYB7\.5<d-5PK9eVGb&g:7VV=N)477/NXJdP(Z9+>7:
F60LLPEbL\RF_6CM0G)I3cXfGcGN66=@XF_a@\Sc:0+4,6)68]_0MB/+O2^c0@/+
X::Y4U8:JTaS[151Fc5G&GR.6W.-CbC].V@;b/E,YWP2O6Dd6#<,gYRd3R8Ia-0X
0@6GYgac>+P@f;(6A-<L4PM;.2g1=GDcAS4^[I@b[HU1MR9C@EGY-7a#MQ05F,Ge
SY_?(#0TeU]8]ZPd7;\;ZZ.dRJ<2@T,D.\LTWVf@LRe64C5K>CF0LBZ8]@ZA3IZV
Y#fG&&SXVK_a^N#TT:PTTVO#dLEJ7f#fH+4CCLORYD,T+KAJI-JZ\\))QEHU++/^
OdXVYO<9CEZ@96bN^SEK<1V+KOSPBR-d3TJZb.aE&Pc.);S)#NL8U,)93BJ5#2E(
2UH53IS5R;1b81^5S)PFX5W+ZU.W4\EME0:K<b<X:f/_V#SC26DN6>?RO#aIBP4S
M-<X9^0I+eR,e6:3&#@,X;U6WLZYN(JU][SF&PKG[)I[3615/A:TffcM_e22&/+(
P:NF_NRS2aAd)O]FHH<e+5@V>VWFf75b_BH=4C;GN7O+DSL[L6gKUMO^NY?5?aO5
Bf1/.egeJGZYG\./#/VS^9U_gL/8YL;_O?6A@>CKM2C@F7E<SRM^Jg:N=UJEDP5P
OP2-#],<<Zd0^JYI7K;57IdMgLS-J?5Y@65d:8=G=A39gQ-<2).gGbFc0#P8C<fg
P[&(9#)\HYgIY6Pd>T^4&/1EDQ\K0+:Qc[SKAKNV)4Q]30LD<X?0\[5b+:UY_-Sb
G378==7K3&[YFXYFEA=Q73PT)M-&J=S]bF(S[+OVD)M51N\ATU>69NH;_=^]3G<c
dA7QAXO&Z0J8<4E43+^CZV.;)?GK5<\TI@eB6@FH68]^^c(#RUN7IMLL@NRLfc55
3J?1Q6/?.O/C8geed)Hd+.1KT].N=Y5[8W9+CTI[BO4N?b;)^U:6,a[OX:/7C;U9
g+[7L.O0@Y1]MUfbcTY:E[g41gR-2ef32YRJ_bE-Td<:a;YCN[3c@:8B)GNeTGFK
:ab,acZ8+DZd=?&THJ/OP,/S7SN2X423O[b/(-:G9BN)KLA74TP#4E4\[--E:AEU
&cEIJ\cS-[DOM(JJCA)S<H?<+M54I&GbSWf_NNY_c[a4HH+UK@MXcB&UM[DNJZ=B
ZA&E@#/a]LG(:IdZHKBFR<#dS0MWg=^S^79E)Q97,_5D;Kc4-4[/_SYJ)[9)-Pb;
-Ee/;X41\_I<@C=[g1_a@0gY0,MQ@g3ecNU>D#)X2_(6HY7_<;YL)TYT:./]A,#)
#KHaX>gRD]>D4gLaF:J>8.K_+>/(?G(DBQEG&bH#QG7AZcY00EFdA9)]Bac>(dGM
SOS,-U0\CD\5R.AJ>B^(A<3[-RMHdYf8B^,cDB:8RG8&]39HHHEM\7YCI.#Q\]H2
,0E[cCFZJ);#)I#Xb.^fB/aL/(E=/;W-0UK#CeUe1GO8AcHG(/6&GbSL,R6<711B
7<(V1D.?FZc?ZMC:2bA<f[JW(OH2)6.A#[UVPa#CX@e9W\APZ])MN[bFO]V9WR,4
,,<O1-Y<XMLV]5+,0bE#HO0cNZ@Fb@)f=59XEYIOc8C)8b;DL;a\He>,585H?L,D
#.Z:/8G.1_2YCY2@F2B5c#VGea;P(J.JP7=.RD6VBOF?-/_Z=ECMYU-@+(4Ub4H+
0MVI<?E,?--?PINR(2NU_[g[^EA)WcO8(3?1XJZ^QY<APPd\<<cFS51A>S8#O8YV
Q^UbCWNJPgGWYa4I^bZ#,9ad,(c?^RP<[FF6#:b(7&@A:/8]K4.T2C-)TOf2#J@:
\FbbcE(D>+HZTO-UM6]S[dBC..K2KIXAG2f.aGF,g)#ELHK\ZN^bOEN/A)?+UA-O
EP&A:E<V8=.JMeQ+/_,+X([[N-TC4caJ-6]P,650[7=:X30^/AAc6B;R.S3dR3TY
G/^8&Kf]N=e4A:DEX333?^He85dI[g4gA/3G)QTd26BXPe6&05=+9:W#XA[G3&NR
a4KTVLQ7]R+/dF7.>6FK&UeKVB)#8Z&OX,3>@DgMI38^XP\S.86S7JCM6E,\:[7<
ZZZ3OXB>MB@Q[UQS\&c>\]K;><FSB&:N+AP6);HD()B.QcCA5.?E]^A#A;^7RCdG
&CZV@<=<-f6E=a2B_NKIb.Ta1T?e4Ld0[eR8;.NN_F[G[^M\#.?eHAO^=_W#N2N?
FLA=[Keage6?RES&eO/3R-_SKcR6Q;JMfLT8/W<NgDC9EYaHe+42ZT@(-^]&<8N0
=Y#^-OG)=F+A&V)8W>[3;b0OV_N&;fZD7;4UT\U\9P=Q1J,752R6/&&[<d)L?__=
B5VPSLObFdK0-JF2]CFKW;)T>KaSKCc>2,OD[d\1N.KWP[:PA;L;0/H.G1fA2OVH
AH?@(@RMVfD;M+fKB0UHO;59Pc<9A+=.,bO=JA/cF)H.+B.JBDMU-).UV]A-.MRI
+SF(;R(>?&Aa?DV9?9D7Y4+,B=/(U6,K.VP?M/Ha\-JEAIOPXO8O5>V4]P^49VLX
V1\X3B6#D1bMVEdKbY#_56(+2V\USW@IWX90c25/#7Wb0^;_B6MW\S=9BB&0@Me[
06CD_U[f(PQ#G)1D8QD-B)G@NO9eP7(+_J\HLafVbLT;1CL/P\,fb551WP/L<HP8
Pe[7[@<;VWYdF_JY&J\.W_B8<\cIIGf,RSZVF.,JCBXO&]]@8a&CC_.]/0&Z\cC/
4cHB13XP/J148,SCa^LcLO=a#F?IB)d2fB9](1EDM1:B.M7[COdMVIJcX+/8c3AZ
7-)7.^3U:/EM8]#?_+WV4_Dc+:@BO@:0#(\V=5&3/GF<7R3-RF:-QA2C7Q.+HTPM
X+@>5SG7.WD)U6FBSZI[T=>LcQB^c1G_[PI;c=R7ggXR_0V25J,Y3LFdSUS]JW/J
PUgZ^5N#-9MT[Y,QQ.:RW+g9;9F-UDI;\fHg;ZaZa;DU8B.^^D[>cT@#SC?(4;+O
UMWUM68a1YOUVWNGY;G.F,0ME>9>aEQUC]Za8RY6V=73\4;Z#,CQ6>48Y8IgGbfJ
T0PI&DHKI[SLW.+;1_)G2Ff=_HKaK<1G;W6P(0;K;1Y78QB1-1-(g^fO21Y)]f,P
a[G^cP6LZK+D-C\OV)-11@&HJe0WFgN-b.4H0,-?/O]R4(SQR#4@^[1Wc(NBU,4Q
01BCOQQGYV,SaR8DNS#H_5-3UIaIP@Y>+H2?UX:X?eLCGUG&/.8TP(aHD(AD8R.[
L,f-9Z(;RdKg6bTdJH,e-D(BC=a]+0K&N1J@3bUT3H7=[.9<Da(-@Wa463ZHV0DE
,6RI:@Q,>CC)HAHM-P7ZLS;6IW>X_?Jb>OO3(52P[67eB[S^_VF]W;T//NU2ELc?
?)YeK=N#/M3K4[a<:1WTd35&ZK+Hf::(HYg7NE;#Q^NeN)-TUPB><_/MVI32VIbL
?OJbd.7.P30Ve2<G:HFR.b3,K5eP@4_.^A.)7-E6S?Y@/b,H(SYHY1DcMa-DgY#L
Ag.G&NQMKZCcN22T0=aD<(6C=)&:8C7SEP+MB5]cFKe@Q.O0:JI05/cRBTC/^dT(
=c@^TeO+f+5#FNcQDJ(7H_9JTP0,8N8Fcbb1H1]S(L2Z4-gdE]dcPI6TcHE.EP8:
G7=3IY52HD]E483(g@-9^6B=^K#0KOeK@fN?0e&=De)-.(2(X\(#(:&e9)\4^@#O
&bebU2@UA,+a2C+7[gQQ>;#:OVUCWV.g<b<W@^<>RQcZ35+>bADUUPPS0DDeC_K@
K8fGS33K4VdRZ;?=;Ze9CdFP,38/4ZL0VI_EYG@+V,UGd#FS252:0G.fH&M]^bDF
HZg5Z]J5EV6V#\IQ5-:b\:GJOI[.3RW<fF9;<V>ONAJG,DT]_0;-;L[Z<4^B-D](
D<T-(8Ge]f]IQ1gVTI/929e@>@BZEW@BXJe3X^f0XNH(9<[fFMM+/XHf;4b>FU3[
23WQ\ZdOU81+^6f;AUg0Pb_4=7S:KZFa_gd<W@PS,WOHb_9edZE9g&1MgM?\\5AT
]&ZE[WX0:/T&(64c/7@cCB(ec:UW79O@0>@A3S?-RWOQ<8J9HZ+PM5UMQb0=Z3;F
?V3<E_YcgU2^:0+CCaM3FQCGUC6&.eLE[1[c@Q#G<()\S1@5W7=&V:D:VTLNIPb.
K&R=K1+BBW:WOE44./g:V0IA0W7O[1c^;#J6KEFYTL\W\=/-J@/5+C=fU(M^5.eK
B]=La?Fdf_1]L@8[RO^e8IBXXD_W9OK#MSQ4/)g(Ub0O&/#7.7d+;TRX2KDNOeWQ
c(7Ecd#OC]S5TA=<dF>XAb_[Q^.,DQJ8.2EG_P@46Af74N867L:J-_UI;0&5#SX6
L6^ARIUUOZ8V:\HXQ#)/],)dQbOKW=C:7&:3Y1X&3[O1+A77GG6XV?M)dJBD@aK[
K:c5X0^8;Kg28HRNF_QLZ#F)agdf[QIEDaB&eWHb4-#?H#0dPT:0OO>@7PN;#T]/
=)76g.;)bSVg@gF4P,aF,2E;7-L&_@B=>]dd1c+#DAE),+#YV41[UBa:IG4WM4(<
<2C&V[f=Bc?)UL[aCadbL&?e@FJUd,^f)6P8V<E_5(dDJS]Iaea,S9>X]S[/>6Te
:UE=>SS1^DY6dEb:U-fB_(YV4DIeSOI0FLL(5[d8^BY;5e^fA,3;Lc(^&N+SM:0+
Ke(F@bPT>L>(7I&3IH(?Q3EagY0c/]\&\ME#a05MOSURcF]#b(Z5e0^)MWObVVVL
V@gHT3XH+87ZTWG^fVFAHZAgI,.4T]+?S7XX9^c&]B<#U>D-4;Od#YJV-U-<K58Z
2Q-c01\Q/<87>=^b=[:FRW<g>FVK\Gf3HE4FCdL4UgAKZ09DOB9Y9W4D,3BX_9f]
K5^5d^C2NAST^6ICBT-X\2VRP@6K?Bf[6;\D&9:#fPD=TPeFGH4:UFGTEc_gUQF4
0BfBHd:ZD2#B:BGVHX]bVaO=WRPS7:(/D4cB,8S0YN-C.H4YK9aLSVPdcZd0(9e8
Dd4@V4C&f04\].2]aJY^A74>V:K9[/^&_GeY1EY<Y7#G>P+d+ZBF02-;R<<1\e/e
HcTd+JUSOJd\84>-+UE_4=G/)9EcO79BMP\-?Y)Z=2^@d9127L[b]fTPB8.&4Y14
3=7Q--cLW1CZV.R/168PXDR7]S9g9Y4PeT=7J4]XK7[1_70H<MT8P0S2&K1=gZ+8
5(7f4W+TNUHbWFc;=ENXaY@?DC>f<M_gQ\^XX/-_T+-6<F-/#aID)YX+#UAKU0A^
7fD,=;7gV5I->.I?U0eUGKY=+b#,FZ1fM4+eLT.UOJRMRPZAFP2TEGa6A-9<[1WI
OA^83fc(fR(J^]/b/3T(Qd)_dZ&2WaHZ,g\Q4F.[=VB\R=&^Z.I7AL-2G/]SKb4D
]BD()4V+BV.RS<C;53XZA7K)3;BKd7XbfM/4(Gg_D-eY;1-2GH^UU:16#>7VP2Ka
_N^DO(GWLWOLAR\QEA#:^+=P]Re:/I-C63P=VZ^gdf82+G+W=@Q?0)FWbe]1=(GO
OY>7fKf)6NJ\+>KK-d5380)3&fP>52K4E)#4O4;a4\H,YR6)=3@F\?L:Wc[16#GL
)_\91I_((Pg[-3(V<U_O3)6V&-T1]<H5YAT8^_1_#C(&)[OgD6?^[]2#=CES3E/,
b)07fAIbO])]MN>U_6)c_QEHI3@2+=E#AXBE&E64[PG=E4T[#Nd3FHDWg,\f_,AI
4cE/P8[e\V\70#6d=DH<3-JdV-TR:;=RbREG:N79\@ZHTTOAS</:VfUFX.LKEPc/
?8KfaIT8XB_+ZeB@[,0g?BZ8R\.GOM[)KP&V=8?FLA/Cc\g?CTeK^PEI;&I^eM9.
bY(<08FA[F(RWR+-1G6A.fE>/ACV&PGS<Pd3@KZMUI2<?Bc]GB14TFV8M@2.S:+8
7R:G)9XJeUeb?/VM/C]MY/c\5D,KBS1X,38NRZ#&XTW1BV)CePRK4gT5.Z-^,H)f
E_XXe_#6:eB<RSc=Z+>5gWdHRc;MXVJ7CgTd&^WG(+Kf(F4QBN1MKccg8;BGWXg@
TEJ,)WFU/I0YbPY(-)<AV499,:d3#[Vd[P[LX#HDUZ3B40AM8)NWdR9(cgQ@83YJ
1<WJc8QC)g+b7MF6N(Z]BGG,cUW-&YM224U4,IfEB]5S#XfFM>\WdNgb9K[^.CJW
I2NF4GU05I0X>JJ\Fb6KD2(P)T)aC8@PYHGfKU[+3a(PO0=BH(?=P)36/Z0[>_b>
f@THTg6&/G4R_(,-98NKHD(EC\b:7RAEgHE9eb<6.f9O0=^3>V>GFTR9HWF9.[U(
PS2Z36?]fD^KOB&,aNV\<c/.T0+AgK43.Y4\9.I@?YgP]>+=FWcT4a,^L-K#ac#T
&50aR0c\0JEJWD3_3?>[60X[DY)bdAM/?:[]3@4+06VHK;UQT(ZCBf]M=PFPDBaW
cc;,KU^.L^8[1=:0&SNd,>WW.MUCca&W:88ab44J-CLeb^ZB<f=<#U+6aH@<Hb&/
C?IRa8Bf[R=G>87XV(JgFM]R0geT9Z2PL6g<)JZG-^P;)3YdOD6;&[^-AY:M>FGO
31/.]\0cP.YTV(0a>0ML)Nd>b/c5+-C-];BCV@B#:5Gg[W;J8N[HAT@7@Z/Edf/-
V^3F0K^gdSKP9<f]0MJ-.;L7c7SKH-BHEVFD-D(]6=D?e-ZWMSc[GND_[CgW@AC\
QQ\SF.GBR;PRCaYcNFfUHCF;X#,1&+6gH#<Q/f#?MFAbC-3C#1Ke#Y7cW)/K15&d
A:;d#)>89gA@M=\0OS_Q?^Q73;0.YZXY@<&VMR0fS)Q6T9PFMU;>[EfTHZIb_RZD
])3Ad6XRaQ>8=4=W&gW4Y@Z(b8OX&A<<f0O<E&CY^-ADf_W/3GQ];.eI.3BSR]JM
G3F(EO?.Y4U,D/)2R(]I1@-Y-@H&=B@=8YZ,+.=<,22A+b3B/B+(77HTAL7XNLTb
LN(AQ-K;BG7G_OJV:\M?Td0RE+D+>Lf.5eeUHQC7R#B=S[0A[cJC[J,&RXLE2QFB
:.1L:K4IOcRETbZ:51V<D,f(&,GEDGR1FEb[6a/<H&+]1>O,-@]cZadE_+TX=BcE
g-C\IB_D-)98P+9X3.W4)71HP2]),bD)5^<@]cc(\FF[7F+-EKF^C=Oe1:,_OZcL
SfN3F=^fKga&I^G(&XLNOf##B&U-<GTX<0fS+cAKTL:][]962OP^X-RBG,.IB[5Q
,=J+<]RREfbG:@]OSbB?AP,8b^]MQ[LYJLG#XA6<GQ>O2/W1PHN>0BXe^>#37[eH
>;MF#DD+cZ4MZT(Y3VNO4&S6Y7@&0GK:Z3f;JIPLa-1@]+;0gH]eD_dBdDb3>PHa
@_H^=1+UOIUGG]a\E]\B-[g5_7ba?+XAN3,2gW3f[H;6dKX_bMBC#QFQC@]5<Ra]
C;2[2cF;-[[7d=-Z=f=ffT@,0H^Tce;P^>;0PdYWI3-_K\RT_.3\a-G1,?1LN1#<
g.edYcfMAY@OZHB0KdNdASgV25Ad&HRQNFWJ)-a?MZCL<UZd>(67^RMHN0/+Adc\
)ZA>d1Q),RR/CWKQJdS5bNBNI^NO2JK1TNO^&[;LgGc1J3e]O\./>1)]dZ\>>O+(
+7YWcAM[)X+&RIY)^1G;R&PMSA@QO#@Q8TM?_V2N.@])(6Z.(,9#;?#g[869B3)I
fLV9(Y@,15DF<,Y5WIN3._e4?MSH9OTf_=1Z/g9S])+^HaQE-#89C[R&5LIe8DA(
)+>D=S.M5AB[/LUXEEU+J6TF59c\2AS;V?AFGY.Yb5V+Q5/H;H>MP@IaYU>5QQ=>
QPOA9(S5[6?Tf6J,3HIX65HVbT&35RC)PQ2=DbD#;7I3KS9=5aAVL)YHeZ<[-QEO
1dUf)FWf&QIIHS4g?D,#M57gObaL.[IFN<YS5GYFEA\Gg7e6;J><FZ9ZI4?N=B@8
gWKBW^T)6_c+c:>fPJdNVX^:5,Q[.2<9^Z31VR]^\?0M3(dJ.];2D=/>R2B@7:HQ
E9X4NgW_)0ZBXHPJ/--/0+OX:9)[V5;AJQAJ=.&CXNOGDW;bLHD:T9^Ae+XWX<a&
Y[JTaS43Lc@IKd\CFC^>>ePI1E,EGACXYY]RODZ-7GPG4D;/8-8Y:OR/,PR/,@c_
&:7HCHR^Q]7f\</XU&Z:_:M2@I]6CfJ9#F1CA2+-MVEH.?D:LRCY18G[Y?/NOQ5<
^KFH61.L:a?_a0_5HM/a/QMKNB-I<?>@Xb2,/UI8/@JQEQaB-U1F6EaVFfIW.<3Z
Xb4G&U](7-GPCFM[I^F7(2Ec3-Z1GcMGVAK8cX0IU6aXbFIQ90I,2.C@.6T7F/E/
-EbO6,O^=^^bc)AN>NcF99-P7aL=B/=M;eQCROgI,e2^b([]_&4d#6IbF#T@1T:H
RQY3Q56S&9S)5V5-#0Y;P^DI]&TF5HGc^e&>.ZGe5V:76dVaDQbZ?WR;/<M?BXRN
&5d?^&.0\S@C0@gG]SPU3QaE#Y)O8-+M:AJ:KVCJI^99L>&]&Gd6T(I^]?_K\OMM
@D8160;0@E=^M/@MUa\Q-HD=AHPag(VVCISd5,>Q<Q/@gUZ06Ia[;J&@da,=K)Ad
a)MJ_@YBTE]PP3B:NO:@c@B@@FRVR]IL#b3^B&YeD&5>JC\Mg?X-,E@W^L&>5GN<
Xa@Tc<^;N;e9EcDg]?,A_V1G>QR8AQJ#AZ&:7DOVC25.-1a34/@_-W&R;d>ONSYZ
BC(&@1A)gd;FPBCH184^b5P+,6G<XL,<FW1@TXH:T1]#eKQ7GQX1NWG^eA,.)22Y
QIHL&U;ATCX2GG;A,e_3c@YA4g,(S6&^SA@?ZLR]\J)<N6^fKX(/T+UULcU8^/8_
HSa,_H=UM(96@RH5]ZOQ\+YYL92)VARMDJ4=0?[9/FW964;[A)>D5>K76e7-/G?S
[IPafEdKHY3^AVg@.EVPW8EaWS[B:dSKcPcZd@5,H1Ja;)P=:f)TW29KPI8MUB@[
_/W;Z]PUNbabFLfF_G01:O<\6,#CPC_IO;U)XNbP?Y@49UG.bU1NYAe(QDO2f_Y>
0CCG15>3SQU1WXC2dO8V3@7aVA^A^\YLG\;agf:>J<#[Ycb=M20>JcTSHPFc?2-T
(9?XbbD+)<PQ5aNN1M,(#;6720Od#+DG]?21K-V0BQUAKM3X)\9,aN^5Q-]/c\.?
AR5XRNFPN]QF49P1<UM[_]SRXX;/4cRK&F5F8Y4&/6FIeCJ0=^7@W<L93NgBRNE7
RKJT3YTVdHN7HTU3S-+;:ZJ4ZE]fS/,JZ#=gKZ1,H:H18MST>EKNCN.>W:05IQE8
OX[Z9UIGQcL^?TT\KN#^E;DAV+MgXc#A;A?FMX14d2Tf[L7.aa:_R1e>L.I8[QMK
NSETPX5Xf)1TFD3gE#9^R(-5^G],Wfa?A=.ICe&/T=BQOBaA.53#9/O+4X2HfE4#
aR?CL>7Cb[X+d5La\B?=[J68RLVA9E.451._#>\>dMU9O8+J&YH:Vb_T/V2;Q_P?
dEA;g5OK>,/=^B5Gdc;:Q4dU0G@CKPQeUN>8bY.UgDg.3-.KI9T^d]^d;5P.PeG+
2EH:C8f)\affaA#f@^?4]?NFZIa)bTE8MdLMYQC,U5eS4_eMf8Q1#^<WV;GTNHZ=
)((3;1D_]3.9fE)G-CHe?:W?6X0XD9[8Q:5\[=Q],b)TVWTZE1<:-8JKNRFW]F8d
7>NVQHfZ_f@B[3\C;.EdZ6Vg+V\/_\B,17PR@YNEJJ,M4d^U0M=-IYU<7909+]^(
E-E>2BbGd)49_6CYb4;&?^ZH+JcAKSKL]IH\cg.J1,VL=\c9]J=4#XcY@DD7MNba
4__>eMb954R<X1U59OC_3f3K/ZdQ84HDa/2?SD#]b8RG2RBN&6T@)f:)3&60UfNE
eG8,NECU40b.4:MV/763U3B,9E9dWJGGCffH8=V,PAdXc1NT^PX-[bbT.6H_W4G8
B.(HW8/1N6]7a(E[d_]AEc0\=^._:0dL>)6Scc2L^&-F]cEfY@Ee_WaY_(WH5Ib?
Z8&8^51fB#TeK?5_f8OSFV=)O@I/&FJcd@FST]Pd1-A@=;=[3b#YX?]8dfX(g6]g
<\dI9?b)C/S4Y.=Wcea<5)X9V&&>3d@6WRb4G+f,PL7=]=6C3]>ZdWEP8e5BX.F+
fSNM[,0AY(9ee<?GVOQ@egdcG4CJUA1FF3e47___SA3KSJ0.TA,;,<,7I9e9C\MV
]NF8JP\>=H-6Y+I)YV:7\M3<Z@3GEcNdE/M4JQST22Y7:>K2#L+>D>]D)K1/WP#I
aYEZ)H\]\F.f=4?]Bd)\]J7.WA1,Ra@G+W@HZAGVH&F0DLE<-\GBZSH>CX^>U-\K
e-+c;#C:[6E\WWWV.OM^/#/PDH^QE<5d..S3gLJ)GJ-=GMNEUffNg]d^GKgZDf8e
JAR?9\I=ZZbQH5\ZgQaH#1(;\13)&?(F,K#9F](ZH1AbU\.cI:5PEXKY:#(7X+0@
_OCaL6,.DZ@Fd_W33X=Jc<.<75E);e7DdL2+P(TKMVI1H9-6^2XDc]c?]XRgAeb\
4^^?Y)U&SFc:ZHC#2?Q(Y0cb&8J25]MH7=TgV+)g_ENcG_P/ABBUBP7NHOG)=Qda
f?+XZRB8,UgAXPO,&X:V)?\0]/DA^O0@RZG##<-9\dV&eN.8ZX#5Ze1:;d?8=A-O
L)WKMdbBJRB(LKJ1]adc#/1=W<\OP7KYSRF,93ACQ2-S=M7Mb(A7fW]WPY-(UO&:
1?]4Ca8c[Q(ECV26L_3#WAG[8E8W52F#3;B>(g[9b-8bfV^V/XN8>7D&G&<bY/Y]
.d-LGQC?I_\L_EDJ9(#.8KbR]<:0?+adDAEGQd.9H+]f5eH70#6R(DG:XKAQ)2BT
Z_KQ:WaV0,NSGLZO>M,ZV4.F\X[R5e(d^>L1,AH\G6SAL<fI_Q<4Bb?@T\V&R9Td
C<9>RaQ-^J@,_;SWQffH#dgTUd)P@9\);\4\ZU+M0=4c&4-Q11e]O:-g(>@(906U
#;g2T,&B&;\PR?U<X:BLfTHaE2\WILVdWT^83WGZcLC&?2<7J20Z@PJ5V^/;M+TA
OPXe)ZEU09#R.??fae@Dd6POC/9&+c-78YLHZQ(68IG<-)_9&V2.IC@]<Sd;HJ-Q
-EA^0GON1;0\UA/6LB8=D)6\05OF6:6C0PH>:D+?,TfVM2f?(E8+U=J]1fP+3CV:
9?W2<IQ67@J[e7&T>V@Xe9ZH(?H):OC2(;f&DaWUMdF4QIQT02B4I/^_=,[=6F]g
+?]Z_QBY8+N:3LOL?&LJ_d^gF3SE7:T(X#X9&5O[(MXRObNgVJUV;SI,WJ&^S/.G
O4@25?7fU0IfS6fbcYePLB9>f.da#P2dTX@\?,J4^(ZB:/4J,5AM)14NGe[[Z[Ge
YZXB)[+JaYPLMaXTS_KX4]6PW;-R/IFX\D6@+Y.&O9[\G^F,Ga^/F4/7;NcLJ5MC
eD(LGMBWd[_=gCYgFPFdW\.K3DP3@ADG7587W<]0^JVWc5@LDf-C[bcT&F5V,3b[
M?4/W7:P=[g1O/eSD-(A:bg7KW<fW_cS-L#\.0AH:/NLVf&gAgc4O4\7L_Xe1X4>
D1;+P.XIFdC;)\Jd,JMa0-?FfQKR)2[,>/T-SbJ=:U/XF?-KDYb2#OeDeQfZQ<De
;+.F]2.(_Y6_<bQ:N<HLOTG&#<Yba=L7]H139Ke.LX2/1g#Q/S([/RQdS#O+UP4\
^SdaJ)#V5=^XW9d7AJW)V+B;497T20LN8E@J[@?VF@V6Pb;W5(8;)\fOC1g[X8dQ
KaPCB;.JL#NTIVbg)T_\V:2@.C0<>?;dAAeUD0bLT98Mb8>+1KC_MfX>Gd6^UQDX
B<L([X_<_Na;CaYS?NAL7FRN>54]^ZJA-,\=gbR_J9U/fV01U[[N2T-,.RZ/UQ+Q
QKVfVNRB]dUB83Kc8N2Q;]TA1H?D5N<E0#0XV2,aA,]\W)MN#\\,?ae4:(bRQ;\\
U)(B5bE#X1T7SZ4#)0P#K1=G;VJ0I;=Xd[?b0FYN7J3QV^I;0<57eW1eKZ]5fG:+
S:.b&aZQT.D?)6-_8OQV\J.O\P/)0]NTb7=Ja4U<&>>D<c<b#EPa?cZ0Ya47E/F5
^,VU0X_dbc_D/:DPYJO:=PDKTBV2H\-,MAXAc[;:\ffYFCHOc#M8W=d7;2:4]0gH
A-)(Q+O[&9XFbX,^SSW[c2TXYeL8JcG)a^]HXBRcR<R+&Y7S#g4:;]A:QAgaaH[V
90?/?GcMHY)>c@DbKGT+,ID:)(=MDZc=]9@DK9>D]S;+#FNO&I+GMUH?IR:@?4U^
aD0Ig7RX,\N)Hg9(:a#TTZRbRR0O4T7W;)#CBS)&<aOY5<+SZR/b2OfY-P5NV+RW
(Ee1fK6(,HO&/7Z)XLHPM?//-H+ROCBT_[M?_dHD,RFgM7f]WOV2c1#Q#d;WLaWd
^3_C:MM4NM1@7#&U,./&,W(Y>KPA,7cdDCZfA\]CW[\MT(L+L=&_Jd9&XG,)U@.(
0+:B@bWIZ1L^/ggY<((&QRf,<3.W#Vf<Y&4=,57ZCIPg&7b5_;QYVL.\;AQ)(8+I
TLL\;)5[+a7_/,ggba=Y<Q^XbfFcWZa>aSe5>NJE&Sf;>_I\/+ZMV&,#2>NK]@6a
1eE3.YR-RP(W4=BN8>5(?:#_:-eGg)P>G_0NE]Cgf_Q1SYO8)T5E&a_b\P<:S.d,
UKW]NU&_A1-G:SCSb=g:9_-9e5+0+B/BR,B3_\ND=,@+41)Sa6Z+S1FV@GgS6+QI
>\_1R45,C(>8g9PG.GFA6-Q]8D;E9d.c)cSbKD2<@N1;5H@6DeL4/W8&4#NfI,\#
)2_Ad>Z^FJB)6<A?Z9QK1/9.6=8_9M-4g0F=73L9M=_C&(d^Sb91;0U)I<Z#A6:#
\-W>8^]&DL=BNd<JI;XHUY+B&LA9XNKa.fa,XR:S:[B2NIOdcXMb<Ya7?6XR,Va>
76F?6V@\cgG?@]Ab(>:<6c>V5.RY8^2\dH1M^#SY[PR4XEYdQ(5I,BMA\PIY/4fE
Z;B::=D9-N6>DdS5Bb?.JY3JLGI3XI2HGYXVB[cC_5S0DJ+I?>-M/VO\I_TZJ/Y@
;5/<bQDAR,UWU#(2L3=SeB)PG12cG9]X-VfYd-^C9&gA6[^-@&5LP^H_LCGUd)/(
a[MZHWM\/-JYgbKSU(PLPdS6&L29/:\Q/+g:8JFPZD7RDE<>D^D(F]d26(=DF\2H
eJKR3CQ3-1A8@HaV^CJ#9V1\Y#EJ.8E:L\,cN_.F-S^ecK_dV?,+_ga^e#@>8768
7ea-U=D1e1f7<EA2-,6Fd__T;cQAZ#Fc2Ae]^gT0__3@ZOV89bc?eSR_P4:fIH+-
9:UBc&XU>;\_g@47cD?-/I#.4d7;T:@BH,,&2_3295G@D013&=T.LZONYG1YN7:9
TF2G36URS1f3F1]a4F78FCI(TP=PU^+<^/5\aQ7YU[BYS-OC_PbafUI#S)[>K(T,
F:YKJ<G-75WG2I.Q#gVbR@R]c^T_]WI?:?MB+X&3U2JL[9YOa\KXGF(2f--+ET0.
F4.gYPLCQ3MJZGSLU<3:55>(\P<1W@1SX^T8M56TKD;1W9+Wf?(;Kd3BT74:T[CH
2-1PWgAfFT9e+;5A,B2c6A\K.bU#C,dYec8M16gQ7Eg@ZO[dBXN=35JHRdAPS#@^
d?E1/?A/T@;@PS9(b1>:\/ON60WX&9NYRM/A+OA7])(S3K0T/[N//JZ@DBKAX?><
c/]L2TT,f@E&,fPUBOMA3@#J=#7EKMR)b?=1&(ON&MVZf/;ZWOY(B<;aT(\/D\Pb
#e]+#2.,cc>@L?ZK3NSdbPQOJG.?+Q?gOU6;2gcS]SK?1/?D(:@HCa5?=aXO,Mg\
3fDQ8S<ZNWJ@051MS@GN-(Bg+:Y<Q3S<(U(EH7R/gb([(GG+1\8.KgMUMB(1,4C#
2_6+6#C#/ZYEAI(RQ[=GTVEN&?^DM0RN0Z,=cW/[VUEP]A[cb]9R:<P)?Z8(I8D)
Y)ZERE1WWBH#7NO/T+,JXe3,H=#HL_ILT&GP?(/:O83>GP=20>+#<A>V,I<#8N:O
:[T[0D-IQC6M:@&F0O6g,QCUH=&SJeX^+R(L)R:Bc;3<Y-XCZfM)GUIGW(XS9H)?
M4RIG@U\d(>#YScSd5bb4YE]3^_c9MF.f=[[=_2Ob8K&0..5Z?13]8YL4Q8C74JA
5:6<&>G2)eRUMM9?gg:I;]U0[c7ZSNB2IOSD8^cQ[P=[\>_8Q+=[FGgA:4>D]<<]
IK1;#1.>H;JNJAfMD5?7#S4eY4Cg[(K+dVTI@)L3IZ1HM:Z?W]D7ZA/:28.8A8bd
-/4a_e1>5VV9T&;J.L_]bSNB[C(-U6YK3B_dCJ:H8DadVb#0SaKZ^cC^e&I_Z7cZ
,/ST,F5H],#L@:#dF/e=K2X9FOOf3/AU2NZ7+U/3)@FVZ^BLS\7(S(ADS#W#Z_=C
YgT#U551S_cbDLe9)LLEKe30_dF&VN\B6SP[&,3P(UC)=RA7BPCaU3Ref.HP[+BZ
b3NB;:c&[GT^cA1/:WBF5.#A_6G4>[<dd6]J-QS,SB(PE6D_5BeUZ4M=DEYWX&::
>?OL)N;:ebc==0KCWg#5BEVcZQcbaKfJVZ.W,7+GgEX2:U?HQ#S-0S]b;39J/6EO
<Y3eY(dC;4QQA9X4=ICgG]])K7ZD,c3T_D9gW/ARdWQ_FY<))D-Z?J.e,-(++6?[
E7c_BP4R_dT3ZC5adQ9@D:0b[1B0CL[cS6VO^O:7Xa2;_dYcRR<#@EUWFO&SUO51
U.1E162QKcT_d)\WASL]B&HNOC_&e?6ANaPG_9_/M>+[YK]L+UZgIRU#gD^Hg<;Q
PK:L+R;Ac[9TSJ1Uc2/V:&L:W;2ZT2GL^E+O;0<\Pg;WeI9JVTV-g:;F/4AED4#,
>eHc5VVd];Uc)5QC1JERB/H4P6#_]S18D:TM1B=OK3a,LI]^+a@I&6,bac;UU_J-
H+f+.2N=(=,4d:&YQd4AP:>5FG.PYG6bdFR6<DE(g][#4NV]T@06PF(F#(BX(;SA
g<TW;4AR4>=>=+5&@X+#Z^]];/2(<.Y@-R3dO_D2:J\I5+<;+G8<OIZd+dcd<HL)
8M/\:D61Z]?=;P&@K.G(.@Q4c?V@@(&JL15BC&2WgbC7(c2C<M+VB>^8#V2b8T:a
M&<=I^e9MBM?IO&<;:;\WW6_GEDFL&WIDS>5]GUgXJBO]1=<]2dT\Rf&1TUJST^0
Z##W,E]VcR\I1+E[:]+HF796EYPQg1:/XJ,c/YZg:ND1AC.g)1KN;cNZEB3#W:OU
/3KT[4d&L2<-VL)0F#5F)B8KPY5Q@^J)K(<#VY?N=e10^P3V3:gF7aEB/.ag<LbU
YbPVOA)CESA.]3gS.^L<)]K22e:WJa+C)7T(/:&Y_.?2A5]EG7H/A/T\T82\ULWL
9CN<IJ2&]VW2c./H5E;LW^A9FR+VQUY2fE:eVSUKF,+6OEEF2eZ09FE(cMOOMWC+
N:P(ACUL>MX+MSMC^OQFDTPH+f,6(:c)Q^=DT;CXee,+.BbTHL0_OQ=&Y:X1CPgP
5f8X&#7eAF:eS89]0@<WTS\VS_g1PG@@_K4<T4?Nb@ZOffIU90KGWV6:]A+c#X7S
3ZA[\]>LLX#H3ICTa>cWJ/[.SNO&e<41WKUH^8ORPWW7cLbY1X24&5S1;]cgc?TO
4.+)Xb3Q6XH()C81Q[22aeWFO)]2BP6S#BBTME@L]R&e];<L<:HR7X&NTMT7H((+
54?Q.9>/38beg23PNM[?D>DBB0<&aF&d/04.8AOKNDLcF@G>e@SJYLFDJ2(5O&DS
JIO?C6<&;2^B\Z;5dLbR:6TV767X6J/e7fAA(#^@G/,(5V_3.<^OSd4(dI(#ZDe7
W>@IV[\RBVB8K2FbcLK7J8+V^[WCT+<)eWfUCba^d.T+I@@W7THgSO)aS]fbf57W
[S_fHeFQc6:?(GZXd]^092CD,/&=Wf6NX9[LKBe^G^#0F]<N^?7dD&EC7(faV,ec
\BVbQ>JD^]BU]-F(&(a8_)N;_VH1?W)JB1V2V0)T,ABGLHcJM;)J#.-C6R&/]Dcb
N\E_8EME-KV9NI>GXAC7+CVG.;F.0cHZPf0V&CM&)..R@AV5DLQ2V^F98JC.T<(/
X,EK^_=a6XOB34ZVB6&cTQWXL8b@:Q^:?N9IUX11CHT_@E1U86W7L]ZOJ,-XX4:(
.>D/O3<#78,]^FN[S][66&O?]\M/Y0<::7G5A8I2=24Q;8-<PA6.2:FaXCGU(R,/
?974,ddFDe,2ZZeK5M>3&R<LEg8aDSCVT_P&4.A8&3SM+=?/g&L;YM?SBWbV]ZHY
](YKNR8XHLS^Jg]gFgN).C\Z;</E-I8TEda0ISYK;@4TD<0\?J\e>9<OB_Z@WW#L
?XRXXC^F7FX19=XZ;Z=WM=,[7N/K5e/HNN)^MX=X2^#2I#RJ[OIaf/beKC8(d)Q^
XG=(X1A9<d+MG@NA;4LPbP^M_.Z^Faa60L8T^<=2I^N;e]T.:bI;83XZ\=b9I_O7
JAAO37HT_^eJ[b_beWB=RRY+O5K^&_@f2@dRT754ESK7cF143P#::G7-H[5.M=b;
_\P^=-9]:8?Y[W5DN?K2\P:<B+0?LQV#(?=5Y=B/6F-^e9B-P_)9/MW;<P>#Wd?@
MUde(R-FBILPd0^7LENS(Jf=KAK;:CN27XWe:7\dOW\2[-J4a+Hd0bIeVI)L3/dO
JLWdP)WAR0f7N6b@FGPO)9F9CWM1S+:&[@aI_EIaa3)J,T&KH(;IZ_K41#XSGbb(
]Q4-(fS24Df:-ICK#K0.;MWcDIC\[0LXe4g:H4G#4gIB3L=ggMW[&8_?I,B;f=&=
-KeD/#DSF+K/gaeNJe2d?_a-0+G:AM)Ca&Y[eSB^.\6DHX>L@RDf:LJRG4]#/a/:
16_]>Z#[SM1NfSC#/bP=5Ng_ED#/Qb=N^e#-U@8HX?:I0,KA>YAK?1H2S1OBZ&OV
a^0&X_d;RNQEa+c^Ua1dBg.2=E52^L6H1^0]cY0]HIDb9LOacVX)?WR5MYOadGM#
B;H<)FM.Da(f3P2]U=_g-]R7N^fT.[VH7dB4Wa_;13.7g)Q-+(L:XRWUVD[a4,bV
(MNCVX[BBZBff/:,HFD<W[)9/?BO;I@K1]>8-)<?^QCF<H@(1f.V-1AfP^CM0-CR
?<IV@YC5#&Va9L<M+T(I12>][c_b&/[FKLYadRLa^NC=X,cBa1Ue76Cc<MN;\)#I
>e:E877bW.T(]1NU]@&WLY=QK3dNH113-[1e@VBU9XK)4#\D8&LXI[P?8DA=L[F-
_K:&BHJ9#NaUU#+J\,E-M4DZ:X;e-Y8KY42S,b:X4]/J2dZ+dT2&HAG4?TWF0BG+
VTc;>S:LX52#fY5cE,-H]8#O@96<.4HA2Z)fS/SKKJf+MG;HL[:@DcRO2##6]#ga
8)).]^W0Y)]7@KQ+[8R.[1+]([CE23S?>fcJ_6Q3OcFG^WEb/P_La-NHBANGcOL<
W6YSR4NT1aT8^;J@D\:+XHI+>XJ(REN-5Lff7a+PQ3,YRV,6UEA<1Bd;7>0,N-3B
8.5E8^6H/&HN:^UWJPG[#GAdIH4O#+@LJ4LCdGF=M,/X+[\JcT&Y^@e,P:+T68cC
RWG:Sg@2U;\P66W&)Fg>3-,,EMR,D?<1Ac+8<?]OD;.B?a;=LgQ&(0)Y8F7T2;M8
/\X==<(eSeS/8Z.3L<c.ES@A6GC+HU=@#IaSX:,8:#WbG.96MDP2?0G(d./a,>3S
/?(WHAV[2I83GHaJ(d_[&Bb.7;2F)>2:/FLOe?L86/^(;4[(@M>9R_+8I<2(+9@.
]]&+]^C9Sa8/SG3dF[@OdY78XVg,6;Je(J>P@e<dZ&K9-KUFV;fWdSYLA[P)>bAc
f2LYd&9G6(S99QKEZJ=Y.K,,R;PHE0WVEK&[ZXY7[F]G6X5UbXQ_BYa?bYb89/2R
IHQDJ6Nf&aLW8+b#[?T2LM..+LD6S:N0HC?A^b[Naf75>.XTTEb?4K(b\<E:O#+J
Gd)56S7=XU_6gNTOAQIc4.T&OD4LV6ACHBBM/)]QeFc54RVGL^JZcOGAC;AS=VdX
95:[^[c+N\&,]2.B6G/1,[OXA8eaIWS-\8B<fZa,H^XB@V+1,B8ABYR#TJWJMJVe
7WaC:PMUCdCEd>6(^J_-:Z6<Ya:AV0.e]T?F]&,X6Gg4D3\R3-PJ2+(X]OfJb(4\
HDZYc\/R2QL3U_e/+0+=d?B&011C[&9\6e[@JAc&,,dY.:6XAT]+T17acdB\SGfd
<Y9Z0.F\QHfEV=bB@RC7L<9KG009_LfU^4)Rg(9=<S,0#=?I[cdX8W5R=KQ#[f)F
a2L)>ASa8[Q8aK]O&C2CKgWX[5C;=PaISe9eMSfdE5UPX<DK_#UF4OL&FJ\_J6.;
8dLbbN;Z3HMaQ2d;GF;#?/<b=^^9?JgT_ZI+Ec8X8G\.[ZYeIX[>OMF/;:FON_0)
.La?^gI[cU>C&]BI758.6<UE/3d.XK(ROT-=7cIR9-8O2\bg3bJ8aCN5L3HSP.O=
]+U7^eU8]:H1)eg/C=2515[]9a-fNVO9PH=I\SC)4DdaVRRNRC,M5K6)9Y[J-W(_
_EDNQUZ_3,[X8Be4ZgbOUN6K+eV/0U>@FO;QMgM#ecYb>AI,(\4G0FODX3N5,VIc
R>1\R3W;2fd&cQOO>R:VLUUV[BGXM6F=KRe+2aVC8YT5\V>2CZKf;[Y,@L37TU07
/e_U]1g-f_O+=LS-HZNHT_H=-,>;K0Z@5EY;N\d8N2&,GV4HI#)+SO=?TUCM,XLS
E;B--\0E&T-gP0&gJKNK_3/6HXfVF.:Mb?QI@)4/NcO1UV&QAAXFZgFL<R-JP9<0
D3\+)/O?X146_BCAS_UaEA^1KTKU,MaI;L>OB+BU1<a2QYd6_cX73/PL,ZJYe3B2
F=O3f_KV9;[fZA]SL&>bc:1;9X>Ig?W-&XJ:+:_YcBLV_0\b<[DZ2c(6Y;[(USIO
1dE[Le;C\/TC2>\L:QWgfG8O#+#<7\(aH&Lf+?C(,AH5f2^V9VC&NVLb:(IA2.>R
Ic3GbO3gfQ,a?)UgB>;V^G1P#F&[8]1F^6(;(e;G]C_W[)-WM&Z.QOPg<6?PNe_K
KM;1Q.b?<:eQAdULH\RdM5;^K8H;,@X/b^N[>J>9NfB)3/F-@Q^8)G/#(b1J#YV#
9R8^J8L@_9/[KX@6YbB>R3^.<Kb>:_4B(&c.Q_OC[?[BHc7NIEL?\64>O.SP1_&-
A9MFI/O>beIAB.C\IAHJ3Q\-LZZ(e@KAe50I@Wfe_Rf8FLSfNM+J+PO.Wc=e?,Bb
g^DHL8D+/<?]_<0>PUY5^EO>3>,@U&.:?ga#3ILN61#[T6\7<VV4]Y9f3eXX&55Q
Gd,=[f7])ZVZ^6:Mg[4W/YYJ=LMRfG:HED.eA)I].1?=>(b6-;bLXZB?C7Z6<142
1),XKYQ,B_?89F9Rg>>]QW/-&_Wd]?e1>dCBX<b40RBfd28O?^W\cKXb(<F/STXC
LO_O+)5L&]WS_VS1g+)bLSQc419#M4W,.XLJ+<.;dX_8G]\IUD=R/UJ)OKda+Qc4
2ZA6@Qb4^I/@FWgL&g1ODAFMeBcI=<6fFGag8SFIdEZ0WO8e165/;]-Ng_UG>A=.
ZJ7.3O?@]Zb_8.(C3Aa?U6f6]VR],3DQ_L]YVW?B_L-cZPQD1BLA-TObgAE6_4[0
;3NFZg>HGA^gGN0<GfL]JLWI+-HH/E6Nce/N12b#LD1e7R;4;[[)0HBFLK^_HQM)
&aKQgG?::]14HR@#/^K34/ZO(=VdV;Y>+W<?,\C+8P;SR3?),?>@&T7/C9T:ZbT/
]fFPHd1I1K#A=&V_8GH1Zb-,WSSCJ(4>,6EX3/f9[^0.[:#?7c-bE6g<b;I@A?GM
[/K\]R+Sg=27PO=42@b&QB;/KN?PSU;EcNEJ;2?g-)+4.A#5U:+WM-9gLK>0Te#T
#c4Ac6CQ^+H7.GL0-;/K+OIXJGJHB]Q_HE1[Gg&:I69K&?M#d6ca&M@OC1ZHT>_-
03X:g7__1Y6M2W4,UE,9+W_YPTS^SB8R[F\(:U_ARU.S;E#a]VIeU>Q7##+[F/&]
gQ^2^,RVCL;W>>LTFESPBF=V\(4W>Xb/0,cR[SK(R_b^56H)g^2=QBZG<(b9BgHJ
8(_D^X[f][VQ;VI9&FSG#CWGC_d8aTB@XXbI2ee5(c5aeCXNdM^^Y(,ALH(2C(Xe
acP8/(Xb[-.]4L+[OZ;/#@TH7<\QKb@BOE#Af=[Ub9&.1:/=,fEHQg,H)PgJ2[U(
,6@V<G)[,J_1Ec>[DM.>Rdg^WSb9f3R918e9,;cXW6,ET5,_fPd7D75A=d-3^5QO
(NI:^8F5.Y3=Xg;@-e//(\\=YG#Q5F_2Y?X<[8N&/+X1>(0(=fI_11PK.YbXMPEV
UF.;X4I8ZP:FR1f8J;CYN6]<BEKBTbeX;eHCZbRO0b/><++5N#?^?</X3?c4BHAX
KJ=Kf9?B<M3H2:VMIV+aRH_eeN@d.N>cb7;IX0CP=;L?QZZ0,T4/_dZR9>G:#gc[
/QU@,ea:_IIT?A)\<10V1IRO@>AH9c\OA9L3[-B:30,Vd/GR5]2:I[2_?SDeHb>H
B,#[.dF].E_J4.8)ZA@;O6;8gf)&<9I@P&80,,Dc//M/5)gUWAC(BCcY^]d;CH+2
+Fcb=Gc+(64g;Q1Q@?Y[Xa]d7JF@IbVHZ@;LM#(50]/WPb8MGc=0E(eSI&_=ZG9R
g^<9bd+_RLC(4P=0B<=6L>D60E:E:G2f13=Q3b-fcXR,+\X/;71^F^WPOc_AB?C&
YYW@(F^,;VbOCGH4E3G@cUa]3c4/WH1F_/\Sdf5>EC8<T8[LYXD5>+AJD3UBe&I3
)=fe4_,2^,D[:FCZ1Y9\^]Q+1.B9+H9TK_65>_YRZQ@O8d>I,_)7[Ag77\;N3af]
0)Ec)7e2c6AX>dO\[1I.Zgc=5+HX-GVS3NOFa+J^W<,O?cg:ca+9SST4UYO\)Ng,
;>G]F7=X<]CW,[M6KI@S2PYC@98<#--:aEeDPP_J.#(-aE=AQ^bc/,5H_f5STfON
GO:I9[]bG/IE@+TM6Uc)B3@:CG6Q@bIOg@I3aIfO,Cc>g]X&@ae/GKJBP^[^<IF+
6K&f6^I]4Y.61.Ng1/XX]MH9@7\M]@-ZHB_fJ\ARFB+JJ0.E8D8gC[1f]A?.=MgV
S>D>#L@GRY0Ug0.GVTS(5E^f_(&.2HO5<5#f8N;P_TZY]Ed[VS_V>M,F3+_XV\&b
]O&?gf/QP141&\Uc>1U](2:PU0?W+Z[F]_O+Z_5W:H2f:LJa3:K_/5P44L]aGMF+
(16b+E6D7CX@&4(:LY([-J,CB+eS1E5b=CCIS.c_b:Q/O2GBe]2aYF)/BVO(MD8/
=e62=TNL8OT0\R[J^M@33_e)cNb,d5=F&e=OfG12E7b;5aOgG\&CdO@^\^.V>H;g
G]#^AXI\7H7F3Y=9,).eXQaZc)NTb2g+]0<CIEO/ge+_AE&aU]a[Va</^2HaH:L,
Ec)JG)?;VD4+1P],<&+<YHL^)O.1P5I=b,:H8?YY8Y2.-eb9;c4^f4ZFHU+VSR-J
gdF5J[XZ,NS\-S&UCc[de_fKC>+eZ,Q6a=DL?f7#)6K.3MF6.9faaaKX/[&#S+TO
QQ54[&B3b1=63PF@2_dTHN[F2d=&]5I6AD+G5HA.Y^MB:._])EDGPVUE6d;^73b\
ZE7<MXf\^6\F457JT?U[,\\FbPW?)+P\__EGUSR=RYHK.OLL\?[(gP1]BQ?9=Rf:
PabR[=;KA,@D>1Jc4#Fb5SfU.&@C6^XI19Me@C^:efa>K@5.;H>-(LgSJeCL&A76
-J.^gHJ[&@_b_1E=NM0)U0+/F(^\b9TfOE9F43\Y1<c&E8ZIbdGS&c;AJH@IBHZR
E)\Y\@^3b6&9cd76GRT.S12RH?9EgOY1;KO(@=\?4aa7HE[8[;M;=-U2D2X^\(dZ
;g8fYd8L.HLaD&OfHMRIad9<8bLAPPJ2C58-=R#83[EWd_W(;8ege=+F4<eEPE\C
W6607Ac1NFI,Re3.N&34B[[X9&8J.:(2FR/Y8f](]<bO?EDRcVD@daUTQQ)[X8[X
W4(]-UR/]<-1NYa[1\7C-d/HP;/_FOE#QKK=A4Y.=L:P(JKd5:9Y=QB4C>-Ja#@M
3QIS#DGV+[XTAG<:b95(c-&M:L)8fYV<ae^FX=)VQXe^AMWR1]4f/)D5#c@5;#Z+
@WRCC8@N0IQV,PX9Z1S?[@09ScfcTd?J[C</JWE[[2<VLc<&-<@K19-0<8?^2cb-
X/e1JAKc&]US79CR#<YE0G(H6E9(gg7:\?=8JIQ97aRY1RM^46Gb_Q+P#,]d?VAX
1S?>D=&QE_HV+C(\EIg;I4a2DddVF(eM47HQ/]X_<ETVEMWUJNFf;dQ&74#KD(Ke
4WBJ2XZ[9Z1+&9XL01W@CPS_B8WS]U@\BGf@KaG;\C)]N>9R^6E0GW;,WJP>K1DO
[XYNCe&)f#e:e<>-M5S:WLga_6:B5>C[-8L3K0JSB1YA&a&d-M2>_YU285<fM=/\
e12bYL,39Z=Q=^T3BgRG\:GGWMP67bQLG31<JGV;,#QDFBC?_BR[;?JH76[eEJa[
QbEV40GZS?g2>>=I=S4>fF5<1[?Q+8U\Ye_>.Z5A&+fTB6@<bOG+0EMVSgQ=:N?B
f_60-]KUT>0f:]Y,E&e^bdQI:C)\,6DYR=>,E^8_G]YL26S4,YDg0;(IJ-JC+->J
ZJQRT(RE<M0^.Z@T.P1cYg36N/=H1X4[LGfb7?4W&^.gBf3QUJ.F9QO#4gCY_a-A
QQ3b(45FPI(&=^,a5F&.I=22ZZ#FA4YTPReY#Ld?d8N7&IaAV+K>2/QM9)c3)#KH
NG.)B=.S,Y:=]T8K1LXB[KC@^Bd?1c3F.WECUGH2dA\OcAU,IW[O+:B4Z2RBF]b^
OCZKJgQ6c#dbP)+G^UY[MTRK96\^5F#X2OM-N\]?2<+@C<=T18Q14E&4JY9^/bB)
daUgdA8K1VD-_2.@,GLN/eZ8g?5;?)PHf7,D)>[)UDP\[>08cfL2gP:)QDG(f1.N
IVM8deT?Gg\8&51f5L#>e&3c+?[QGEFHCd0YQ_],YW\75@]@5WFSeI)C_:56d2;J
#4[<Cg^ND>g:TMS5eP6I3/4K>@-D]Id39a5N12/WJCG/dCXT#KX@_V]C\F0;2W4T
:8)CAB/^:4_?:(FB392fYHH5fWC=R;Gb?2AdE1U9Z.:fJ3E&H9edMG:,0@84QLYM
11WX,c9[<6Re?0P0(e0CdL\IAeB3(RWdLRN<G]_<IRT9RMYg/6>WZ/WT=AKN>SDS
K4OcO2geT2PV4L_9>)T/(<R@e)H\Z+3d=3=9P@C^+M=&(-M?E)g-7LG1-D&FcTH=
=^ZJ+f2LHU9:Ee-U@0Se)2\WZJ\^+DHP6Q^)B;,4??G^XK)0B/L7?93>2KT5L:IS
UD[@>TRAAe[0R>=-_(dFEg55;f9_E0/I7cBT?XWdOJ,d[50DOL98JBJ0.Q5E=Ce]
A7Q24.OWVPZS6X-F3J:>/d;fICAJC216&g]&;.&W##_E1Z+,(ASVODF0:\?\&eRX
XP&=SH?1)[Y/LZ.-K^#R.ZDCG8IN]APZ#5Ubd_:_R[<@DXVg],1W7O:WLg^c8,FL
I,KPX=;EK[N[E.BC]b_.@^ZNLPU06-B<660P_)&/1bMBE/gWOP.>7__Xe=ecR)Z7
&EUfN&\&<gQ#ZAI9bMW^R2_6g\5?BBNb=L?R4[Q(2;FT6b]9g1eB0T-\3Kbf^McA
MZU_Z67VefF3U&5e,Q;g4TW?c&?1-;=[?C]99#M^U5Q2;+(:M>08B]]3_A/H0A@Z
ASOE71=NI;fD-YN-b_AVRM<:b?,)[:U,c[)+B33S=Z95Te&6S2@WW)6XQ)5=U,;?
I8OdY3]QdfHR0^],//(,\NEEH\b5=Je/VeKC:PG)4/=/DFD68_XGgWB()bJZ[GL<
c#Z+SI4g44UQNaLITS,g)D(0NNK0LbW.#<H00Y:&)(FEV&)-(T[DKDMA@2gX#TXg
YW;+Wf?L7.R8P[b6g8\eeV@M@[^WdVR+CSA&TXVNOaRK]2,7abQW<W;>0-KTD(P[
SZ?ORO[=Z\8:-Q>\:?c>:]=>cg)O(?T4KWXc=e&.R16(+V4Z@0.Z#gU=?g;6U1)>
QC]#Xg2IOc6>+Y+5V=X06V&9<CO@JLR22@\O6g0R@69?G[8VOY.S7S:E1G&600Y(
\8]AZ/73bBc1U.:FK=SJ):/J:/)+927+Yc;(7GGT9_=a;F,PGC3K7[4[7R7EbWDK
[:6DIL_VCfBK2IZ?Ha>]=G\O+6gTK6c,Z5M&I3<L.CQ5#b2RXV2)<-Q;<0b(?H#U
;E.Q179LgZ;/UY;R[YYW29YM9<B:,YRAB<Q.^]]8C0M\13ULZ/53T<[VaO,IJF/U
PGIZ0Z/0K-[KcKFFdH,]FaJd3S1RHLS<be?.K(^AJ[#JL,.0KB/+00#JLP/6#;,)
L<?,&>R98XTA8c;WBYJL@A1/?;MUK)CX:UF3+NHBJ:a-gYD([2aE9SfF1J9N)<@H
,U8=HY7A;@\635BINQHJ-PcH&CP_A3cI(_@5:&M)+=6/a#JV(#/_RT4Rd;g:2]?e
RKcc(]G[?6.=@;8LZ-aF-CT@VUW<PQ_39)/\(QSab);2&^T_U^OcRg\6@3-:<G(>
;E^?efL1^7(^&Y]5Y1gC@2.EF;KTGIPY:6728ZcN<9>0F5gg46Qf3KC=(4[Q;0Og
XN__(0AI/EL3OHPe\B8,78W.)cM.1#gC,-.J2U<FPL+Lg5NDgMW@+73ecO9Q-bd>
c\06@\/(S]GJU=f+2G?&GU^[\d;G=RFA<Je&4Z.;=:FaIb0GdESVOL=<1.W&RA_?
6Ta=Sa>+P2^[N:@XT[_H6\Jfcg.1dg3K8)[WLQWAE@I:RISDZ+UbX,8O92JNd&\>
[dV)3P]O=LDU<D0^-F)&_VT/1N,(RFOfHA\XVZg9.7K>L4Ld4?aUD-/DQ\e.HY4-
(=BA?d<L].8#27BRM2-11c&<?BHb^:#G1O=EM,cBRV?@GMgK[69R8gXf^B-\#1<B
(V1g+GW4;)<d?31A&RJ;;,D^(M?Z\&AC89_>UDQ?[gS?/-I@GV9?>C#@[WOK(,9;
aKf<MHg9J([0bJ:3NU;-K:KCF@W79&Jc)/JO2-QL9IO&5[9);a/@YMGe;_#,=9[-
ZO?H4XNSa\SU?f19,B@>/B5TfK9\--dgFb453=WYVK7E:d:T0CUY@,]dOYZYN&B=
E@IQ5Bd[ZOPQ4=c+BF;ICY35LY/)+8)2b=+Af8RdXb+aYN0F9<eDfNAe2:8O520]
>\P\YJc+@e=I;gQU3:^M=E=gZSR8\<3V9D(aQJ&3+8ZQH?A<8?WW@,[U@X.2OaB8
g8)g@EH@G#N-)EZTI=](,J?L3X+/\:\R8OT-X),;:_DSC:VdU)gaG<>Z677QHg-T
=5\;5F[M(S2Q4J@8)dJW)3fDASMdV>G+dF[XD4O0dc88]S<O.N2M?4J1<]-4_;W=
/bK.+E\Ua1\)\:6A.KE_V-&fE@U/XG_>R?B3JSdU[g]V,KGY,_eOZ\WOg019,I.]
+=N3M47cR_WQ9P)-6ZDL)gaQb2TFKW9CH:Y_1ZeUO6>[\eP2EdOU@gMM3&0PS509
NFa0.+O60b+g<2MZX1\7]3Y02W2M9P0CaX>=KUWcOcWE=S,5>&NK08WE3.B&KUN_
JSdf^RUH]PW708(18HFaZ?.NQB&D4KTEBSMET9eFI5DI>4^N,AS-Wbc8CNdd0OGT
]P<>:.L9Mb_C:M/0>:?+Bg;IT@@:a.L;\e6,PGO@[=2+[GYG?J7-?a[][Ta>GN?-
E@F<?;I\6T1]U71)b_ecFGNFd.ffKAP#KXI)LU?.D9P.I8eLQCKB1&K1I&-1F.gD
FU4:/..1L2-^4d:.c7D)__g>T;WIK+6P7_FMJbWK6DW<=A8>C[[2XQ]O2VO:>d)f
WY.VgZ](IG0S_J0L#BFOgW:cT<UP7g2/<)GT_@>V(4VBf^^3ceRY7NW-aJA2Be=.
FZZ\LfPTNUS/MfE/:B77T<L9<-N353XNNYD[ULc8_:cXE?QH&e\59\9GP0TJa#Ag
MQH@B+.+0&I6+HNB;3269:NR?5+B>AfX0Y\ZXBVUIb[5<C/X\af8P0/LT_^^Ig;:
DSNg]AJ+][Y10++WG/a8ES+9URc_g1ZH;YK36F\9dFM[K5K0EbE8R);cL8:b^W-M
ZPD):WPX/GBabFbZI;PDFfBBd16X4BPdX6[bH=ed.-BW>X0N&QG,+WMbH95H,McL
P+?D#6O?ZPBOQJTB?\OR[(.[TI34;BdB\(GTCW&TND>Ae#f1O#V7,XOMCe.X2LR/
XIeUJdA#)K_&a/^25&@&H?&^TWGLO2?MRK(Q:_@NcX<@25,d.=@3Pd_XNQ>4]HcB
I0.1P/X<-1/;X9\^\@AB7Ja/^VgT9:,31IN]5I2PUY772.d,4b4aA-B_K:TP[&._
&BJ-V=.3N/^6A^A]/GU]c,R4UITCSUZfg)9fJeJPBD@2S.=5,YMNT,AVHaJMMP[=
@RZJ8a:B]&eWH&-OZ;0HQ0,H(V#N,3;BX<NU^Rdb[7ABAd4AWIP^O<ggG\/Q^XZa
8^HO@DRc\b;\2HP2\<@A-?D9QS1WdJg=>a,OHHKA2&d-X=NDSM7Hb>QE?DOGW54_
74NUR7L>#IHV2+Z:+d[[ZV5-;WO;<K<-^KWGOIZ^<-aZH?YM0+>ZcH;>Y0C5>ePC
/_-4QW;eZfZ&K6OSY2_DOc6@J>YR4F_?J7DEJgU[@.J&g@fN6ddH_RPZ5PHe:P,N
b4.ZLJ7NPgR)e<MZ@(I9\KU7,2B9__.B^PRVZ6AD(5O]62HZPgDC1@f[CQJKaH4T
B7A0>K5PUHW3_[=?_K5TBQ)QL(bWGc\bJ]Y--1BO6#4&?C.2D#V@gQb,f<^1JPSO
_G<?A,Y/,ObcH?dF]2G?3[Wc_7XX__eU/B+d.L.&1eT7,-ZFYN8AQK@;Jb4)@<)V
:G]H;LE_W:#bC+4DQ9d8\9N67bH,&&e3GQ_]LUXSdAFb;96.]EG]L082L:OE0e;R
-8?@E[_WcKfQ[)V?[]W)Z9J80SQ-SJU5]VdF39\QGN0Eg8X8ULa]e&)]?&b[)aF5
(Y&GG.]A#I\6FZL1I+^HS1F@7KPAe^<Xd?_bdA1FH1^<BA1]@dVa1;HD3:7-CHA=
^@:=,_M5XFLW5[^E9,_QR+>PN)\BRfO=[NSdd1-X\E\BZ4b(]e<e/E&)8>Z31)J:
c+IW_]B,^Z1K86YCb6)#a^7CLU9\CRW/8#&e,-f#^KTQ]MSa]UND[ec;ZA8::>15
ba(YV+E+eT-=bZ5LYU5FN29S]4#13IME)E4Y\d>]F6[SI606]E1CO#9g<LK5eTdP
UTW9_B;LRGY=3M@[47,@FP]d_5X)ZMC2fO,BLV52/f8..N2(34bGX5QLOUQJcL\Z
5N[&RYGA>&^BNPZ_,UAf[=9+QPW@L^^J[3TMY5S;0S\MgdR+GRF\d?A-L<g]&<B6
W205H^53_M@\?)@0b-?=aF6VX-W/6SCO+DE8>FN,WZC;G;:#8^A<_XY.8e;BH7a.
F-_KcGXB>Dc1M3H.+BB^9&9c(,bg)=70&Eg5d\GI0fMTE>>YBf\/#DFZB(M>9P6#
bF?<d@N)B2G=JHO_2:VfH\H5:8>Z#NA8^TU>@e,[21aU9(P+BAM5cR]?R;@57GB(
AQ/516LcO&JF6C,Z7#\ST/N<;.Hb))94HJb(LC4F=.Qe^gOUJZ9H^Ya@;C#g22T]
&-A]J<4KeE1d?/5MY/4YXEMb2J@C#:542P43aH,1=NFU/#1SNGa\Re-)&J(108,>
5/Q?RZ-8K@,87R#_\#(/L=Ef(dEQJ32[4[bAHV6W+2^MIF1-g+4T3S++#Xd&@bfX
4]W^+;EJDaP,VM-NEWM,99_PLXYEB]/WHEe2LCc5,7G+>UQVK:P8;:05Z]a)[Vcf
H,\dae/cfLCWL5\EB#>=G)>G<eF&Ze^F;OEX^E.,[PP-?DA)6_W/VNA@^>d_3<Ad
,SOEf;,C2I/eK7RE>e1;b.,Wa9W+NTL_#O-6dc7T)3,WQEP+O_IM^PN9&R0U-6GF
TaZ=,(JZO)5^N#7?&gKe^Y][XRDA7HOb+NMc3GIRNKMCEG?JY1RX7fTIG#T9L,&,
S]I6M\_9WWP_D0T1H(#B:J-MRR_?S_QJ+ZM)-@R5_8L=770#aB5[.(2.^7U7+J;V
^dHJ;U\F^DNM^V05O/e>@c,6H)2K7FIMQdg8BeUWg.T>HBZMXDR@F7OO3KM[);HA
[QfG4^-6/KAMW?##fFZd:1^a0VQN>YG@]TeC1I<:A9&+)^J]e.J[QcGcfG+#L6Y5
M,2.Vea+(<HNQ<f6O);#afYd=,X+[,\8]9@7LdaN0EEDbNPRF:(Ue7M-W=5^_)24
Y?E_PfP]K]P?2<<b.Zg87Sg@8DXc-(EW2VJ9(0N6M6,;2)9+1S/>F@K)S(Ie(/?-
e7KA1?/8#?#eG^\1)XU5Y=a];f5TZ3B?P_I9&(?O9KO5C8eDabNcO-/1M@)HQ[0b
cF<(H:LL==<)&4C4fVaPR+Qe3SKO:YB@[^FGCN&&#XVDZ=T^/QP6BFVe-B.<Q87e
4Q1RfBbM(<RZT(#9f5A_Z6_IA]/2,K#e=QBg:MH6eS8EPd[@P:V?a7c.0+MfISbH
Lb<MH;VJ)<@9)VN2FQ.=G8RCFV^Y;>NF&TV[Na;MPa\AEW0;b]Y140gI4,9#1@7I
S#V(TJ1RR^a-a:HXBG/:AbON2[cea1c1BCY,:>&XcO9YLg[/SgB(>/XVeT53=8)9
ZMeO^9.&]]c7?2A,]N6UKM6,@803P[CLFH#=FI6=H1Z6M0Z>T_R^K=.N3&I.:4\S
;TVd9EAa6HeCA8U?8DT3H(;1LX1[Nb66Y[_CXK=fPALKZbaM)>P_&Vf6024U@;2P
&4I-K)_L2g+7_KJPb>G3bL[>aa(G).O@7^P>_XIFY3ESJA@38_W_./VbbB?da&f+
AAAOQR;d],0R^1YMfg0SfE9fH.I+8-?N3O/9\;Ef2eM=O7&4&^B:#\NMK^,XD?3L
7QfeF+2##KI-bf9JU[&HIN:O)\V_(Nce4cG4;a)A<.caa0GZg[2X;g6<LN[IOLcC
W+8g1-S84NK5A<3;>fGI/)d)#.NRb;>O6<XQHE]H<Ce6_T\CP9V3QB+IZFB/c4EX
:YO3<:,F=?=f7UXNBAa7aWP?9?18,V55FZKT;gKN59(1W3>^(-D;AN5IN)]=a_<Y
G<RX9T+f[bRF=e^XJ+RB7d<Y+S.]U@-be5&2EE0CG1]/X&>=POVIVF))R#RF@2GZ
e?GBZ3;AM(B8FB2^60PG82<91HgP[2T6XeC^N[J2,b__B88V<?QU:;VK\9ZPN[N[
=gQ2H6a&<2+93(F._-&H&e.Vb4VgMZ?.:)N=:DV[AI?#4?SD48IRgQ;[8T;Z-_R?
O6(<[2RG(N#BEN[BaLa#X9,;&2C_QV95TE0ZVFf]aD,1g^F-F@CQBLe5<:^L]Hg,
=-&&\888#F8UM9V>PD+QJO,NFF)NadAVHLLJ:R38Q=Xb4;;\,YRR;6+d\0Z=\W92
9?@gT<+KXUbG493S[9,c\O=LPb6F7)#d^e:?I0G9>Q<a;Q80bQ:?MP4d;VAY60AX
#[XIQV5<_\?W9bS>E_R^4PZcTGRP&HPC<^[5Gb6LXcGR?7<JEP]2fg=3.bC[<:K6
0QV;J9bgEHXH43dIg>^Jd[1SS;+f@:<8f>YI#a7(F,7V4<=6X^d7LF&[1Z=(R\Wa
-OUa<:/36=L+\J4I#c:eaKd]eXUa/ZD]T1?_KLKL=+I)7,2,&FH8S2aeI&8d=/J+
A:7KKcVWEE^gAA-aYO/(2Fe_O?WX><cK+[;,HO;Nf;QN/Re-3_&;&R4;]gV[O\aI
]b_B:?+ggM1Z&9_\<R)Q(/E0XVT[2Wg&^(0&WRMEb^E<E.B)E,(XEN4A/(>?B(Qb
@Na_(QMfT2+)2R2=\QdQ]W<&b)>LOd/aOC;33:US4c0.b+.;Cf8\-,fQOZ.A0<)W
+FT;3d>:D/SF?^NRL\&.1;)eC(N84\e;gd9HNE;H;WGC#I8H+#.YT][a)AZ8.3CP
XK6Ac/aUJ#59S15R+YGMdZAg^K4PWQ18]41K\FY^2H#]C]c>6X;e]P>QI6Z-58KT
/Y3?ceB&LX1>g12M(eF@4dSQ2RKI04B:+U2Pb#>5f>+^7ffaGV.C/\X=JLb71U&Z
P5ZNYbfM]WPM?3)A7A.]\EGDN-dT@=QMN?HNd:@1/UX0VY;.RT?]g_&g(;YV6f4f
S,TZ<Q<:B4B4RTT5Q(^=Jb?H=LH]]Y)Od;:^;/\_)QK=eBddc1-KW2Q0Ka:]7ZBe
>N9Y:9&M:.85+cMGA8@17)ZN>LTU]CC@9J:O>^Y0#P_##U#LU_gOXa+-#eYc8HRQ
L?&LeA33:7g4Rb?(QFT7I-3?EZ>NCV(R5dW#Kg[)a[T\N>8@NY:F;.(^=I-_a2XK
8?QZ@U>9>FXba7\WBe3/<[T,J8>-e_ET-G#?)[I]dCQ)7LEdJG9A32)9B#++SdH1
0J@/dGL&1F&aJI6-e&/]A9;5;I+:TB9D_/DA[V9e]:WB,6HLZR\_.Y[Vd,@+>Z09
[I+NUIJEY/>\4Z.&F2&gDfHW@:,[@=[HHaCS+Z>/69QY/.HN>a,WY4f+^T.D)<CB
GS0KHRg8+7+LV+@6bTOXK@X057CW(A;UEY5XF\ZU^a9G>\a/G>>5II:@J(C/780V
I5X^8,C._Z/bNV>=)J83=_#=J[IBY6>#DJWI(U;@JUGag4_R:5O]/1X\9?T^AbKS
c2JHcA)_]77R&9.UCE]R<dLR^P-ZNZ6,0#/\5;>X>>7/ZZOda#bFZC(L,Q(H;:48
Y^7?@Y]8=M&;GZ3]>Rd_(@-LLKKNbGLUeX),Sf.d0XDH)bdcBV.+:I1=L&HJ8[L2
8HE@TG+U_Df@-<WO<.?>;6[<f6Td>fg\@/5KZSL77_7f/[ON^<S_fN^9QLZR^_a=
+N+F#5>1_&IV-MB,(gA,@fA1,.24eHY\OXS]KT=SVc)<3@Gg[+D9g\ZO@:X6,E#0
#2aCLgaWJ=^EKJ)-a2\cP?>fIbNNQPBWa\6cg&=^<c8]U#B)=MV#?8@bdPGZSGFK
0GgFfD[8BIM5SFEgcD7\.6eVV,#C1&[+^_@4XIGY[=?_.Hf9d).0T#]3W_gM;<3+
HK,LcYb#-2SO^<4[0\8ZH5C]N-?[(/G>4e;LV1K#7G44^Sfd\@51dc4NZb3E])]X
GS?eO;82^09YU-S\1B]8(A/2]TN=e/O(2UQ+(:&=F1^ffQ#(.@Fe@LZ:3\3.Z(E6
>eWD2,H2:I86WATM1-FXK6/6K1eH=LU]IYAgY10GgX2FC8[.[O,XG^/40<F5=6aW
=CAQD/Z[SgG;<Fd6_1J@)NN.2D.:^P@\Ra=Q2C1]R3aMOYf;LC0D12B/N5:Bb^SQ
cFK0,bRW?B66YT6>FOGTY+ZJf6;^]4GG-/(gBcaNfUgF3GCZ)Z(<>a6,d.e;+<e:
>d.20YX?+bR@XLSX+c7BT>K_2@V)YCW)RKT64a8>b&KOb#3/:8?d]g)[RV:aMKQ^
gIB/,T]JTAeW9RLL6e^YWT;E68@g:d_4:W6,BLgRPB)6FM81c=4UMBI>.3WY;:[N
TZA>[;\c:1b=53V9,COK[KB2092:TKgZV?>F([_EQB(J>7-+DZ)LdZTF02RE8PM7
-ed0HCI\,8SfAILgD\]JX[eJV-;I]MON:Ja@GZJ_)5[,Z2gTAa+Kff8O\8OA&4Ha
D_F\6)dR-C.NDRg(GSS0.F)5ZN5@.](WCgQaR>7[9dPIR0XC0-,PHTHJ>USY#)[J
P4953JO7P]Q[-T[@O+RGYT#TN6SOfgJ<O3;#E:1TTb8PeTDWN)(VK_ALC6UN0L7^
).;C8#^20/_9#c(#Z/\+9d>CfJ;0f1WLX=&RAMFE;I4&f7D_Bg<7D[=D;D3397G^
>V?EgS.1L(>2:=,71#O[+ALM<Y6V2f;T)_bD2M2TSfE1bJ:U]Tf:3C39-Y>OUM8;
8(3]+WG.D<N_JLe.@FAO6SZIXY2e:D]e+?HH^09CbIeYUD+JH@.X2B4F>CV\,X9c
A9U+QBCV^+8&)D@)K9I?5#9G?B7OE-ZdR,DE5U)7^+<.)_<&OW.PNI9P)bQJa&Ae
&AFNG4M>LL>#G0=IXIGMYE5@LH0(?,W@[LUEJ&@FTZHJ.-SN6X@0;8S7MM+F7bS@
)M6(Y5OgI3b[ZL4L0gPB,\-:2@GJWbL(]=4IPD.CSYIb_L(H_@S2#H4PYWWO4,[4
JB=7f;:/P85e4I@8T;PD+P+/<(b0+#WA5gGP7.bK-6<HEI:FQSdJ(6Ig2+MD&32[
Vc\PHK298/\U)@:]#7FGFHMZ:HPeI>H>64?<8\\#5bJ)7gNKG2_UIUg>[TOQ5,YD
N##5950GKU<Dc[@V&\X,;6JTbT2+2BODUD#.X@?A@QB@U-b(^b?YP0L),0C8:^@2
_51NAM@W#XL8gHAa@8,(9;XMR&9),bIAfgUE##>R]^e43HVfON&YY;15R#OYdJ3V
Icd\+,/318aAXT^)R9B@)>IY^<[2F<C#YM&<.41#R/AQ=8_;HWGf>FgJ+^-&dX<^
YY9\84ad:./X]DMW[(,?U6/\CIKEWYABH;[-FHI=)8NFC77ab6A\@&2W,(7(-:,8
3).O-eV;MPNRDPA<,9;+3.g)?[<eNIbWRc/#9KM_a=SVf[D,&NP_eAD]3:=Ea,YU
WW=a1,gV.8@K:?36#G]H8_7?J1]<2WgC5Y]g32DXI;0fB,5VNSB7.49gdb0(^QJ<
agbcga2TP6g_E>?U(W03C2H2g5PS(:XRCW]:290O[Tdd5]3MOS(AM6NF#f@2H:A1
_\-SL?Q3>#9_[cCEAEN=L]>ZdS7+I<60dD84<RIA:>RGZGF5-GQ^U(&2JZ&,a97c
RU_bC6.^ZAEb-&#K,G?G/2PPRaCPQFCd^e/aE6Ve?Y(I&fI/:0g5ED7R+@+7T_R8
Xc,>f_J)=_CPF9a2HO?c#&[I;+=PRL&7HT^)P4,^d86UNU2<M]=J05d5P)1RFS#D
I@Hf[&J#_/34339M7#Zc[6OL/;A+95#fFFLC<_J(3f@.EZ@WRH#T=7I\Rc.+VM,Q
,Fg1F+F53-Le9TNE9D\049H(_JP8_a&Q;4&\XWZUK@8Z9XMA_e4f^.RKbI&-dP95
=P2BdY-6Bf6BbC\9L2NT_>>[S)[(9IZZ)aPUgDgQ\).#Ub^V]RFZ2/H^\I]L7c.Y
V#eD-L-&S:4B<DHJ+BR7/NXXf1>OfD7^gKg;B8R^=aXB_X1f9Cb3&g3]=;D-;&a3
+YD9.4ffYe9F(@7f\?G>a#HG)eF>+L:JIIC](:[8_WDR/&E[.7WPC@CA<\:KB0a/
<[c7#DD+Xa\SP+>7UO&3][Z52B_BHJ0Je:LA5[&SaE]<LW@^g1fa:X<E8cEKBAa9
\_/c<X:.aJ#RP5dB0_OB\dY@eERS87R].\LNKBHHB)a]VHYLD+LR^+.1F?a323.f
BX47]0<8:Z;I3+S;M4-SVBDI#MAH9]5S^EgO=5361>B]a.5?B@:=IQYB8Yd\/Q.A
fEWF:]c]HIFP-?c&KGdgF2.WfLRZ(41c7Z/HFJZCFc5Yb7I[[RWF#=<WLI-fGS5_
OF:1e55SUO7A<ecO)P,@1K_&UZe:>^7c\HLW]c3]aY)ZQT1K&LY38+WXd^AS>A..
Ua^,Pg/G(J5<4?MfM\3d)F+9=Y<NMEKMgd29,R>A[&UAJ\43PX[H0KM=(Wbc-?\g
<9GQ6EHUNWQGf,Mg?X[SRdCM53]D<F[ALaH+36J4.EW1,eR7Jf1^XT[BCa9DS:+L
>N()/=YW38gLRI/O.+.LQ(R,@EM)K,UaOXZcZ/[DJSE.99IR-T7bBYY]e@T)EBP_
[eNZU],aBM)W82A6AHEN-Y>DZ==JD,953DW+;2G+O2@^^3?c&cMEX41L:_?1]T9-
M7<,C;E47+K:H62c.,FC+@F;^Ya0C,EFW.HZF0E(E.DCg]aIH\Da+?[^GX.PS>(+
0GeBA-[<W1NU.]0DaD.g+GHU&4?A5U@-&#8:ZH<[C0<^/dXX4Ue>AV\Y<FRY<f0g
928L0Jg(g75;1f82(3YOb:7HR9(5N1\E&9O=_\=>=bPgN.,VF<\N1c2A.MB:8Oga
aCdfKeK@KQL7IKdKEG);FJ3,8Wd7F;)6.#VB<9584NF3CIfER/&.KT1Kg/g,GAf<
8g;NXZW=SM9_A_2+E11_9&[QZS@ZM0C?B5/DcYK2e\O1-(VFVNcBFYN]L):Kf5)P
3J(;_(#f<<?B7d>&,QXO3AI/>7&UC[Z=WFT:KCVI2TWdV3G7@-89(_,ACcGaH;fA
_\7-FfP=NQULG]9>J.g=^Q8<[D^dY,E\D)AT7R7X^,42[MOR0S00T25DR@gFP/J7
eH,3DIQ5G/fE4:KO9YIRD1DFIMQU##^&DNBY<VZO[W-gEGd0TB[3M#YOaZc;g<A;
A4)#D/?;6^Fa,dH/UN&=D@(^Va8W@VeEQCI_1W.URXg8V2;[(9T9PMC;F=7TFC]e
DbC3GJ=7]P/#&67M44L..13ggOTHaC0Vg#9aJ2?;:>V18-_^a\YbZc;>ceMZOJ\O
TeWfa-ZXT-^ACFV.AOZ,8^8[Ab-P_.=7Ng+&)17X9>bGP1cAH9.WDB<TAP)^ZO&_
9H:b_.[+A7\U,eH&O+9KODT27d7/6MF5F]4WO5\SFddZ,=IHe4W_Q[JZB=B]\,@e
3N<>e,OD(<:SK=19AU79@ECLCf?6b(HW,2/TQK>5ILUW=#=_U?0Z(9ab=U@[X\K^
]-+5GS3925_e7=.&??_^b0<PdA:G4B6Ob+(2=3]+>PGRZ^VRQ1I(SH8Q=[+1fED=
H+d@bE;Pe<2DCIUZ(dOH>HbXKY279GJW3[Ug2JY[<eVV+RDNL2]G\MP=N9,+C]Gf
8F-f?F2b_Ze3LcGXCY>XE.I3_7EABZ?.>6#3\Ac&c#(I9WH=Mcg;[)e8Ddg=QA4[
A03^+X[fMVB_Q3H(gW@C@B1-S]>O8)_[X857EM9@?#VAF+T9GF?L#E7&38,GJD:(
0+A5TX726gaPOF_>Q[+=3g7S-WIGPTF1SFb,^J9M_;cBNY,6-P=L;D[T=3K[O06Y
UVYgK2)B_BT\2MA.eK0OX1XV?AE=^RESeY]1MUZ26;HLN1_&,Qc/bY,&feIS74UG
D#=IPZcPFgW3)ZS0(g2-/Ag[)W]dFX-c3g)>TJe>==d5:,_Ge3>R+e(<_dPVY_^2
4eOeVTNBN0Hf8MSR)ZYH>:Q)]=a8#L+O/NMcK\^&H)f2\;<Z10^,4[O^OYg&aLP2
-a=dL.fM=5&3BJI(/f&-8#:_0992TbM#OBae>:I+;8AJZ2M</;a@8=B)J9S?^(<\
<g\XV,T2S0.AO>=cTd-=B>H)C_gEg6e^L4:cWSe[5+O3?a5g,,25ga25MA/5Q5T^
(_/?a5@PBf<<U]ZP?4fD0>QWFL[dQH_.TWSLU2aSDKHUV)EbSR8FTU,:^8YER1B3
fQbV>K4Y1>SL,MVQc.FQS2?7:IJ)RE:P^#d2Z\[_Y,5=5?S-4FRaH2+@;Zf+ZbJS
,#^SGWG+RE0V.Y2&4Qfg9O)N^#HJ6(K>Y_-NefT\YgA&)TdL>Z:UWINc43(dS-Q4
JTI=#ZCQaf)eUf_=1.Z3M;Q6>D12,8(K70YQ>@S/e6SX@[WHNA7V/@-gJ0JJU\bC
(RMfeK?TA;c/M9ANE6g0;<FcD-IeeZQH(3.Gf2)LZ_UATM3I3R;e+63g4AX^KGP2
P5<,KgTL6VgKL5HgA-&>HcJF=,N7+gHd:cMY]@=4#beCddT=eQHe3\SDLUW@;9^6
F>,6HXNVT;.]>I/ZbBe2Xg6G--[>1b+>5M6Ub)(7Q.#Q:gb1KJWI8/)Y=\HZ^;/6
1PZQ]CgA#8M&11VE0bW^>A/OM.3.1b.O-DPae/Y[@56gSY6+>@71RRI;AK=Rb)3>
XUNSO1YMLWUe]6><gGgT>g-K5O&OG9dQaXM4KH(bRAKYC\,V8:b:]3^P7^@EJN^-
I61LXZa;XcYD&N5X9N5GTA;.WU@0W^5U.[fWA-&2&OB]A>,=:SZOU.F-+OVdHe0]
/9HR:e1VgK7@[^ASG9BfX;L][8Rb70Z_L_E=7,5T&NZZVCMPd]/eaAIG.]Q.YPJ=
R/U2BNbEQ^&7S:.b[UNV3>N@82][V+,6Of;Y,\36f&U])cbPN&fZ4X7P41a[E#R3
,F#B\?.XcC^U4_\L/NN\).(C;@PQG:F-[RLYMcF0I>XOR3603TY]L\26J_2gb\WY
S8&V>_VS6C1-5.\d4^R&:/7:]Hc[E_adDb<g<Z=ODZW2OHJ/LG60[]I<6UDfDD9g
g61NMYfT8,3UcVWIY/A_1(D,f:S>D372FB8Udg2?TALR)b[(W=H)X-+NTgP1C2\P
JK7M6b+da9>@6[-2/\N\SRV-)=94F/P_1Z)UM_E9Y,TJ?=/ENYM?<;VH(7<Y+RP?
-E570K&L_Zda#Q+Z4JA^6<.]:caPUMdVefWVNCYOO/)CBN0U7(D475BKWIQd6^LB
@2J1;FYT(FNS1?Wc9(]\HXPP>4U^b147([6ffLV<6M=gW8SME/7,-?0?a)@=_add
Q5@_GL(O&_K=,A@X>7?;G45^Z1]K2(0[;^edB58#&^U2=?L?R#f[0Q8YZ4=?]5L,
4#=><KOL.4&&0bc(1gS_8.NRE(#>5XJdP.\X&CNUc)V6_I#W+K1]Dcab5<5O8(aA
dEcWf18#=Wb9V:XC>=ZNe1T;1;-ZN.&M^>I/[-d=0WB4D+X8>fEEG:#6[;19WK7#
VAa)c,5Qb;EW)MZ@-Y;8^0Ag:?I31Y.e2Z_V8RR\\4-5\5CZO:9AI])3U6VcE)YS
=/:5[K?DSeM##K87Y4SYeA<#]a&5-YRFEOdPg;b2cA7_gD]G8cEcB4/,D:^]b_.^
&OEXaY[0GD#_eERYLZN^-R07)F[VW@4[CfEO?6F)-GML#YP\PQA6,J2XY-MOIH+4
>cJQ1f=8bCg=EWf?8K).\RUBD#E47&T<KT+?+GFgG:D-[3/I[FU-C)<f5d/gBd[#
\,GZe:<#d>)A5)B-cS53:;HbFJ;IL4bgK5PN&/HQM2O-@,T(>11I5[YC@fK)]a?\
A4@N[]eE3b)FSYcZL>BGOTAX)[[/SA?(f(HF(]-8Ve+7KbSN[CGT)QGCOg/VYX8V
IB29PQ&-XC-ZfbVZE6cNO&3GYfMWH66SHfB70aZROOf;U0b[GLF?5;U)JFaRCI6f
5<YRdN]D#LPV;-I+0L[FL67JQH-:9a=OW^[&T[KBUJ.C9<]8VGW.C\gPWe5(7=7)
;cc.eCAC]J[<WASMYBTWRH8<gFYOQR47g;\eOg)()PZX\X?-gZ8H6Z)NAQX;-[+_
-_).J<G\YO.SY5W+EJgUfBWS^-CK0L\WD\^5^&LQgUNb=U/BCFL:6(;)8WC<;R:9
g)6NT#D)=NCg2(U:a,2CJV9O/=C2F+,U7LEB@5+\Y<Yg2c]113IMMBCcL\MG&-X@
J(_K-[PY6[FbKbC=EEf/e#_1bC<ZC?]A8K9UUH:@WOBf?++-;Yf<O(SF+bBaeYF4
N@Kca+;FXR/cZ@@(fP40RURa<EN/<BHK?-cYM9UcFJAN547e&geZ+b@d--5G_NgB
^.e>74g3<W(/1XY4aO(JDS:&@fS=]]^Jf_80PL],<F>#GY>HWUCC0<:)O0M5PNJ.
c;(V/\J]^IX=4G^6bb,@OZJ;.,ESY_D#IIOCMM/E.bV^E5;)gP3]feN:+XUYNYV,
dgaTO:6cY7M:EgV-L7][RFDHIJ:&9;23O5F7]R-UL<+eXSL)#MbNFV1.C-R9_BT&
S\Y>C&.G)]=5[eP^@)[+^_\JE0>QZ@RLABYCGY16c:3c:)g3]J;e>\+KF1TLP(-K
G=<F7;WV)OLeF>AJHbD-L2?&O?ZPWb-=+;2bN-[6.\YeJD_bIT<1MEZCT4+K-GQE
R\Z]+bIO)=@cYVJ-De8YeBXR.\B<\P6,2Q)cA3dP4<SHVUP/R]\P]XCH\c3:f#[1
1PMf#=e:).(D\?HW.+CHVA5dec9?784[U?/WH3,<e.8f5C5[>[XCf.BWda\6(I7<
TI.aA-3K5GKE2FM1[gX_L_4\U9IbcC(]WG=GQ+U>6DY0V)K?^fag-2I9ENBa3VOX
OX0g,]GK16AgII7Ed\b\g6]D#PEKL,07NNJ-;3L9T7Rbe(1dPQO;f=@N+[FUEc0Y
4U3Af8I4/3^UN0MKUCgI^5BNGR-2ZNc-9@e-?\cKW].OMU+N:dVX5.8@J]NgMVTe
R7\IaDP><5=CG_[@?XLbD:TRY.JO(>X2=/>ZfYcXQM_TCBU74aYfDPb#92-H]6_Q
gEd81[Z1[<D/@(Sb,\+9&8_9dLU@)/-Z;T4<E-8fG3P[]AZfbE&D:e3)cAHNHF]M
AFBCWMY?cE6UL;(K;AR[W(JCafV/>d?D2U]DCYP]5KGY&eWO]41R#TeeX3-S_Oc#
F9T6V=Y2826D;fS;7WL\;&M.@[#_LW#_a3^:6=]@G.[g1fXS<Of^MgE@g/1RN:4N
D2-a8[RVJ2HIK/6G-LHUU=8<^&<UbFd:WM;R-(Y]ZDcUK#?GR-2+W3?>VW]KWE.V
V7:&P83bVU_<RZY0^<62V:14JO4I>#TLK.3AW5:WR:)D>,__9#+(dg>+BaVIRL\G
.^.8Bg-@K-5DTR]OUR3[d9bC#XAGLJ)L@&+e8ME?7e=>g6171]SGG[XH8K.bT@DC
)5@P4?(_/LXYYbU[U]25a>?#P+WdC0H.Reb9abae0HJMbFMb5L;0D[>Y+ZX]L\Cg
Z-Y17LaXX.D:#2YY&Q,Te@P4IY8QBU3fB/&a./dSDb-#EO1LCaKU?+c+3fDIC8dB
-9/LJU6F\_HA+-:SG#0&2b^8K.BSSF];L,3&3Md_TWG86P.SSdJJ#LO3IK\\@0A1
EAH?(67#dP;L3((cNDN?20HUB87\>QeX_BZ>3Q@P2TXNVQD#QbB?JX9)=PKWb<fD
d(f3bf6L_O>4=L\\5EQX7]JP?7&JL=VFad/)e=3C3Wd68F3/_&8gTQ=L5=g8GKc9
7:,BP)\dLc@T2F)<)URO;GN/<#<^-RM70fET)FQ7DBQA)GWd.\+If:.V8gW])^X,
9(O,bgJ(e&7)A.SR>:&ZVf:CR8]1:@Q:/\1M45gNdV^?XZIPSTZZW?+f?YN_O8I&
c7^gAAfMJT;_,X)<\=BN]?PQKKU[,cQTa-5Z0,SaLb6d7E@5&S<=<E0NG6T?X.\:
db/<HODd:^^O[KS&aL0c_QT/4L^[,/LPY8.BH<:2YY6#-1S/b9&\9U3^7XK+3ga,
,Z2-H8(=8OZY.4NaF<#N&CBY=aH-fIDAH&;#(\@WT^&K7;EYK_YP.-TLIBLg^?VA
<fM227:P\-_1bd?UgYW#0OgX=KAQ?8+C/&20I^9V)/;49#bD)dXC3MaOXa#&aF3[
0B]IC@2C2]KaX)[(Xe1&6AAc;9U[-3F.^NI5&6Q\&WU:9e5ETR482JYSPRdQ^Ab>
,@/CC+JTC,3+9d.DdLZZ-27.N1,&60P)^bg4g(.OX/]A?<Rge9GWHQ,,(6Se#U=O
FeLcWd3dCcDABUZ,da^a^a;6ZV[_0I-(Z)d1cXUC;871WcCc&T&_84d(C&W7b6RW
+V>36UMG^86V#]1X@96IPN(#+@MA.:4;Q<DQX\c#?FRJEJWEW]g:ET)C9/,VM+;S
.&N#PY8Lffa#Ed(^G7]-_2RF#<3Y0_P)X(Q>1T@@dd6#D&<>1.+Y--6.+4Ob?OY(
+7BacS[BLfgU+ND\eUHKASQPP0MAg2<FMaX^YRVeAL3@Q,QK1/\U[GJQ3He;d.)2
b?]9(KO5Mg_/?;dAC6afWQ.1=X^VDdKGEYP6/034YKF?UcJ9A_e-Q.:F^bDL/aAK
e?T+.E9N-1B/@/XS\[F0EH^Jc@DY=T?[1Q-/VB,aP_bYS@[+Z=,N@+J?J,H5U2SW
11ULF7aB8TJ^g+M9KU0A>dW#NKVD;I:\G_(dB+^@+)0(g0P/MN#?eF7bMDJV>WFW
=@G?UMK-R,GQeg8T#Q06<=L^ID=[PR&]QEY;W(/O/YZ6WV=JV)KQQMa,_2HVQ2I(
2f>3bd;2-1>gdJPdI;7@ZML,U[Lb&5]b4OU1KAE&K>MR_(_9OIY33QZ3/PPN\)5]
THQO\<@GL)fU)H60RTLWO;LU6eQ#YGg\5283<V(V:f_ZKIfOJg<W&XFg<^A6e<<.
Q^F\[d43U]_NgV:L9;+<YIeGRC]&<(C3WYO/TGAEPILZ_/;X:=:_P:Gb<<>U0ee[
_aL9&>e0bEA1W>QH_ZZM8B):_gPV/R?E8S&E).K[G[[[T7HfBM067SN?@Z)]dII+
D#9;J[>JXVO@[a>b1PD?=dU((H&NDbT8I2DKH0?0:Z=JUM8V?bWeV?X5.Q\@K,=H
,Xd]XaS]CFca##3=N6^eC91.KKeFI7]]]6QaJ,6QFV4BX-5a-e=B7KK+c+R;,/4&
0/704W>C1ANV_UWZ)NIBgff41J:,KV^]T\SM^44?+ad)56R=CAYSNUPd8LOQ(bLH
#Z5Ia.VS?0cNBS9BFK?BSP[K\(,,>[6-T2K<?[]fFSON7bL6TD0D+I6KIT>:ceZ5
P?b<TV([Z?eNE&EZIX]J-@(CF@.AWLb?Ae>bN]UBJ76AB#PB.:II0eEadN<T(/I\
4D#9Z__H[&EJ^&T7Y1:aYK,C+9D+BdLZ?XE+8eK<;+TRgHJ#YZF3cG@W9F?bN#+4
L&g?C@a&IXT;(d;T6,Z<N0#V0,9<ecTU8?b2dPF3WK0P>#HR[&M.UD7X@)=9Q\Z\
=Q?#YA@IIcDa;BUaD6c8T)1aK@eSJ0&VMKHIQ5:PbX2ZaY^1,^B1/A\<X4<(KM,7
50PB9BOD0L]Q5D(;<VOPRRE8#78RHZAd<-W#75^QE082DRB]+A]8D^-9Z?J6L(f_
YLgZ4ccW8fJJ@5VK>&EX7dCPR+NR;,b&4^c]ZQeHKQ4D+fL9TW95B;9))d2VFY>E
XIA7;f^^7V5T02@RS\<RfA;gSYJ/O(3L1G37TU,Pf,bBXDKN0dH;Z:8X?V4VW@+D
0e=FY(WUTH1K5fD:Ue3K8<\1]0UE]&#D051g,<N-,M9/.\970.3T)R\.@aVEcY(]
LTHcKH\26?&TeA+N0BC95[JG.9BCbQCB060b\PF,F(f(YNV?Z3NAG1^Yb;8D3+^b
9TLHUHfB?fKVST0H]D^g+e?2eM1>;U@8ecMf487AIKW&PO]]],&:@5S[?>GY8deN
c?W35LG)65F))8eT&73:9O#]GD_3S9S2Xg_?.g-_(1Lb]CY7^V,O?;^\(,.)\,EK
G??<6;0L8V.-#CIeME8:_G(N4JT=L8f(T6Va-VAAT1<L95V=]-XfNZD3\QWG2:_6
L^U\Rg@0[53X99c[8T0&MXN9K&3(&fM=_[+WSF:f4]?<K6dVT/1/>K9JQ5AAcYNU
G)_>YR1QJU)\MT0FQ,LAYLH+7>Z/4JH(AS-G&0J9NFJ0WF6^7=G@Z@PR?Q@F:b4\
J00DP=aRX^U5E;.\W5YZOYKON);\I@U.42=YQF&6e1@--0g.MO_J6/b]^<LL22=Y
+B;U:K8ZG;A,e\OMRV5N8DFHFRJJZ(0K>A@)-cZeaTCb,8PAU?P5b(M;F?Q_E+VN
\TF._DJ:aVV4[-\R)0ATNZE3MVg?U.(eQUa1^LV)#X0@B_CG#LWSgUg/fEb2_#C3
A<QV+QKA0g2V-BX\?IKG31.+4@6b-#8bF=-A.2]Z0M;A=N/JW,4e@2E.DJ9TVB#:
D:NY^F^E^80Te?7.BHJ,](X-3BUF,1]QJA^G9V,:S[3TYZ4,-85H[GQdPAK4<-0d
VIZ+4D@1HaMJBPGgGfSdQ<?HeGMXE>f4&+@\aIdB6IQAN:DA[,dHY3^&N[TVH8Af
->&T(TUCb7)K5c8?ST:\fCI9-[-K@4;>6<<8+LVN&T,&QM2SaZT3B;B#6bf<BG]L
.N#f>Y9QbggV+ag6GXeLE2XZ&OW^29[F<F3_+I<EeNdC.((e\X_#a=?d:Mf@;E?T
>&)7(Q/X5,B9TCA29C>XX,W7BE&aA9Hd0gD5T9U/H.SEcd^9VH&&W1:[_PZPVEJ7
/5HdfRDgQbbX)<TgSQ;FP&U9.FIR4dUOE):;gc3-g:GJGRG0X.cgFTU[UHXNY_8R
V4U8Y_PTYPKf#D)#fR1:Df#D_==&M9gMbJ0fZ=CC\0C:dG_<O,L1INCT&.1N&MS5
NR2)fHLUG>;K:)&@?Pf+:7e67V=(T0)=>([X#G6fDbTf8SM+Z:[]QF)bVRU5;9^<
KEL_NZM9gC(.N8XC=<a9;,Xf:-51A#[S?TVPO^f(=);R)I7W=]_XY9WM&ENUTC8b
]7fMf;EKReH0(b7(<ZV+:_K>=6MCAS-JOcWL3VLa3V^HF/QaJGDN6INI24PW(&B>
1^PRC#58(,#g(AR63f./C(]Ff8R7TJCE+]NM^(VDba=4d)LRC)dc70Lg)7-XQe0C
K@2,b880LZQI7YZK>RP+E<&Q\IYDBID+\aM>b(#6RM^[@KV6e;&0Vb3D>HW&RbW>
1?_OL7Kc@\/bI0L^@^8K@(;Y7e7YUIAAU159:F_SRUg93[?&dFT#N?\<B4&ZJFLD
BebZb/9CL7)WX_HGUOC3dMS3g/+^cUK>a@@<-^C^bM\HC9U-=C/&<IF8N7/2CS>O
9NMM7E=D;-#BP[7(T\^OUYfH63Q3.5P-cL@Nb-56gfXb,DIKeP2G0Aa1_C5SAeSD
deU&2MU1E\C#6L4=:aC-N[OY\bP^a3M9ABMc/0b+\MR;IZO=:S:4@#;J./YcX?&W
c0aaWFH920H-V_SC)g#S7G<H>BbO]:++VD<T?4&2;P9>>=(5JNUZ=1>S<fY.[ea;
VD2J,>>DV;[><)Q.0=515R_GP&.:4JgZSC79O-C9(,D<JbC0B68-#c]S#.@[8[DW
+>VCS:Zc?LX]-4I.a5=Hc-9_=6G^E=1,)Wd]a_>Yf0C4E2CQTaBP&16LV0Ng(_]C
N=H[?)P\\E4>:IEg\a\K@S@IegISd7;S8,WN[_^&Z6#6c:?0PX6[^RcDD/BFQCg?
+fO/KN[ZJF,R@<P:b],;1TZ_GLFQ]RUF<2f920(Of/?-DL@1f\N1?_8B)P^/3-M9
G+=ZG0@1VZJ.F_C.4&9WKZGC^QLJB=9RX:I\g))O+eKU::Y7O;b(+_DM--C&gaS<
D_NR31W(a&5K&Q(88_A>O)(7BEGX]UR[69WT:;)8cS;R#<,C6B_ND6KaaGU;JP+=
=cQ5LPd__DF^_^KLbJ[]&2;N&^H7PQ?T)LFZ3?\a0#N@^;/VU+g4[,5-E0,@VR/+
3U[F-Z+4UD(NX:3;;I//@0XATN^3P+P+[KWGbES1SZ0??1.gcV0>F:e=?\);813W
Te<7\\V<_<RYB6d+K75\PXfJ?,WgZ-&5#=UY\KZ3V94=/))K;=O]1[G.<BCC78=K
:K#PaBJRC348]?.eCTO3^4=U=_Q>L.6Nd9+CDYd[bG\1g4a-\[B3D;.M#2R>PH8&
c#N9T:MEcF&SS-T=1G;<dHOgd&bNN3-WBHcH)A_af9YXfc)P2U:KOFTf8a0:COQD
b>ZR6]0NF1Ja)E12T[+(?ZQaF\H<W09YI_I[WbGBYZ6J;I0P6(\U<W@NS7+V:8BI
QG-DD1W-O<#a734ZGD@<@Q?::)aUZ.eLUCRWd>]PdY.2gG>?fX:>XQ36I0;0g_0M
AHC7(R69f:&X2(1aRSQ02)@VJ&Aa3VWX:ASYWOV7G#.:.4&Z<b.A?84GAbK?[P^N
-aH>d_?M#>/aJU8GNSbb/NUeY\[<b([3F0^BHWERb+):^\E9WRA/HfLE92#J3P#B
&Z4-F2@IXF3=<5/aCV1\8ce]39@G?[JB[^/fH<T&3?1NKE+IFG2J/FJb<b#S7CY9
eGY_7E&&/\5aQ8Db4A=T(M0fL_ZM#Og<&;G__LbdB?HfH8^I\Gg]3\Td4FfBU]=L
\A-/H<PRN)e6NGR#117VOZ;VgEQ#=be7C@OegMV97+BSC)LF\JDFLa1^gO9OMgP;
1V-I9VJ>I/7/W1PZI:0F]Q)P+HQOC,J-?e27EJ>TZZ3QaD=1>TY]KFbb&U3XW(-)
6PFg97ag(A?.20.^MO.\f;:5gT91BD3K[VLY\DR3+00&]Z+B=EFg\F3?B(S+3_.b
e2a94<YGQ\X?/dCSI\[M)7:BN@de@bFH_DTPLTWU+F[Y:@W1R;fd,-g,J<DS]SAd
<5FM6)CC.-(AP(;J96Y\#dHE=_OeKOb=a;G[S?:g&ceaM)D(e@A[cV(GD.F5Le4\
NCP)3C98R?bab_3?#<Q)OA^,T/d3M)D[^T,_TU\E)D=:,HQgM?Q_1PR+31:JAF_O
&):4(=5A24@PVLO/#9<?BN6+/;JL<fT:ESgAO)a3&_<RL;f,/4W>Tc?8>e8EW(8e
TUEE4df#,C1<Y;?-U,5C+B?U<8aS,CU[Igg/9dC5MC<,Fd25WJ)-Ya[SZdS:?U>^
MfXC&/UQU)IAYfFdIK3+g?8.00DSd,/#]WCS>N:DMOR>bANVM6L>[df[G]57a7c]
F(Xf(+(F?]>fM+6@8MS&SPSZ=6UPY;CE[EGGF0Xb,WE)Y<b\H5D3a;QRG+VFWV6\
S?E1-aQE)3HEF]()R:[XSe>1eSVRMY:72bRXd@KO@NQ=]da0bR[3+IDT;9OAO]2L
)c=?H5Wa1YdH#\.W\_KM7;PJ6gA2?]>VfV-X^4V?5Yb-ZHNO(NT./PKH4]C4&(Q1
BJ/4&_bHH.^7/\dGJRCA6O\+a>XVgcH@?cc@=_O<L7Q_JOBEb=Y?PI>MTL-(9NS@
P=WQ;@Z0C)HCZ^K3;(D7DZ]&:Wa[^2=MGTV&d&21&V6@Sd\>1D\HZ>IIX-/2HaT2
g(Z(+KVcRM6VD@eX_RU^-<:VB]XS@I\&dXb(UP/YRY:EFJ,^)=MQLKH>P.+DH:(:
=6-(Df5^13.@XR?79-\1)8XR(RUa>IXN6BF]b(<(FZ0C6/#QYAN3<?;_I_V>Yfb9
7aR.KYe30,YV=:.FLeIFd_+[MKg,bI.3)I1T@bHg8U.[]WZeDLD;W.Q&QY\A.b[d
d8A.Q5HUa3[U8DD?UB,>&U-41N^@R:_(@CF&??@8<QN)].UeX#I^U+<<d8=Zf=+-
HfV#_bV3#a<95dULCWW\<XEI&[=M=:@UOg<P.Y&PA7AHe1Z]>Eb^D<ZCX1GYZ&N:
:<KN_2IA<B;P<\Hdb><M(]VXdWG4fDB0VCQM13,H\#J[.K\Nc\]KE;X3dCU[(UWN
1728<XM\_MIZMc[d+D.QJ)M1&>=Bf[]b1MSV9^=I9@\K=ALCI@b[YR+X9YX,+C+[
40T1IN[Ib>>S]^0(&Ugg@<1W9BR;<=C::@#.57A#EE-&3?2HP>:@957.+-@gAP:J
?g[&&^a^=5K-+N<YMI_cW1>(bg3D38?SbQ9TYWa&c@B)4+SS9XGTGN:\O?/a0I(1
d:08fDccUH_fHB>c.YO?&&C5<2,eb@AfWHCE&g[1QYW/V]+>_\Z,)I(M<&gO9:Y<
0?S5,&6#gX\(IQ.OgHQGDaMd:BB\&Ra^J+#_@#e2?KXQU:@(S+X+J#5SSb7/PGaf
,YE6WbA1U-A6?[0#<f0X29>I(1\Z83BdQC6&.^.LFY0\V97(\;R8910I.YP]X,0]
4f;2(H?^GQ3HgV1Ggd\<cV>:0_e>P8;41]8A2Q-9G[;M5a?<XJLC\Me;T\bJN\]&
I_Q<@?[IET,B?9EAcUVc07U9EgC/=gWWNO[d;d>).V=_aOA@K-]/73I;YFUU/8bA
^5NbbD\7([fT(B0BWDBMJZ3Kf-6QK^O@+BN0;IJ-bfObCCUH0SWO;:YRa>>RKbNL
D-:g=8+FU^E2Y;MReH:Da&AC.\9JE8d-O4PfS<@,6#5UK;5;8B;D.)</L4NX0:U3
]U]=cI7W<;GQ\68^5VGb<bYRSX#aHEVg@:0GSCd0@2M^R2+f830JZdIb(VW2AdNK
?33ILa2,WR(3fZ^GTeKM+.[PbYIH\8e?GYW&5R]2,<H[-3V(Q&^c?6CFTAX7.\KO
@[?JW6YS=F>U_#?8A\+Ue])Vd<=\B\@A))_S281-Xb]3S?HLQ+^#&&<:+Se5]173
0NO]\g9C7DbO8XOb)VUKObJI9\RLY?>_dB=:V7ZEe:Kb^.fc\fQ-(agTV.80TFFa
2=#1dU&[194MRHe^+I(a3@FZ7=bBg9?-I71&>DL<-^PA\ccYN1D@/.YbS7_FABaM
@SW)MN<[](E(O7)7e]S1F[HdH3X1[]+GU91&X)-?GC;99eGGdYSGO=H,\^f\DaIf
cP.QWDUVWZWAd6>5LB_K64I<J54LG9B@&4[IN2O]ggK_N\SHHE?,(M#.XU=0Pe3A
G@Vf5S]?<R::V6IL@)R<FRg26W4A+Cb;T)TDTC#HZ:SecFLXA/CgEES1;WI+AH<3
;)0UW0KdbD>,:[BT:]U?J>4-K\UF/cQBX<]O7[N^gF9b[(1ETJgDQAbT=7bE[DS?
/&9.>O,MfP^+X3L^YYH6f,X2_7@6+34^5/N<[4?\^^O2OGCf:8cX1dbS3CE(9bWN
I(E)LPK@YdS_&R[=50H0>LQIG^357-gJIRdP.967<ZbY_5UKPd-7aB&-X=.7E>_f
c24cNKdZUY^g=f=]#/:c=5B.DV10LJTT#\_A^=29,cB4A+cV_XAF(b76=P.FMI6Z
J5>Q7^H]eHA6S[B3]=(SEcDNfb)G\2_EA(79gV0>eAY>T?Q6S57YEDCfg>[Q.dVd
?T2U?J=ccCC=T^3>=@3;J\4DT?N\U#Q?I@4_#2.ITKNU/\OHSL0GCQd9cJDa,HQB
@95W_WdbQ\YI+Td887+YS8XdWb(F.ZgZZ.bM&+#-9A/gb-U^\7gE8(N29RLE-+]@
+?\K&[=/#@2;d<OXP9KE62,7K^c,dLS6##AgS_4DJ5NW?OM(A-(/E<<1=VH#?/bJ
.I6V>^c8+=Lfg3D#6M0/7Q\=NQf1SI32XGQ0RKS7CJNdI>Y0CO>B9EV31JHWA]OS
A[@_c[H;I5J0^bC.fH#@P7B;N3;b5X_FJW.?L,)X2d]2\&R=<Wf@:[[WO5^02dI9
PEWPL8&VEQUWJe^V)[:C_5+-U0/XW4Y#Z/0:6-D?C9fZ=E#VDMM1L\^OL:#DbA?3
_@]WYe@Y<7)Cd5)D+S=acaY+&2[R5;ZD8<:9fW0P,Y.ISRb60M\8@(>6Kd2)VVe8
e6S2^J-EB]1YZ&W,@Ae=0MTcb=V=I,8((9]UZ@@XDMT4[?g(EGDR588?IfNI1@^<
ad:Z]R+D&:NE[fL(D7V3)7,_&M6TE(@Rg6&/DAR64/N^Q[68W/1bT@O6)a(H>DRX
HSF[PY-)f/(6?c9MFd3CcIe:M?g4_8PB0dJ?Ib^\X6ac]a/Z=CTLfN8YYSGK3Ha#
H=P=-XR_=_D8JW>g=8M)ETfgT>6+M1MUM4JM(5Ld[VQJM;5_DY2@?I).R6(V-[E.
,-[6WUGN_Q1\D+TKDc5bgQ1cK:cEF&#G,MMN?fKCKe0fNdLE__8ed<H>ff4N&-4<
/()MfceDFbTK,-L(6YUb)2;O-^=E^M&/30BT;^9UN-6,97@.,03AY=+eH6V^]VI@
We7AI,0O@1,HBb0>&eaU5b4(=>;eNME]P)3P9gB\&;faIgN-_3^fAg&(UOggbJ)K
]BP79Q+7UYa4@-I=9XOBHO02JMDO\7P1F2\bPY.<[2#PI7G#>JFGG4NTUb2#U>,b
:LVL@38ICAK.bd^6I+<Z?L<.^@24FYAcc<J?2>09/W@[3<0;]ES=7@IQfXR+S4PG
eY-^XUVIU=V-+<H1ZW6S__N&a^3UQe:63G+eII-.6=4\]W^#O3[e-11)0fR4_X?S
DR18P4OUGJL#5:0FW6bO,U[cQ-N8eC3+\=@MegM:OP7U&838B&Q#e0WccO?^Q3db
&bB#L01B@M(QW@IM^eU_ZQ<XH&0YSPF[e5dSQ^[7.601)gHYM+b360YTeIIY@JLL
.,B,6b)#eNR/@4P#B6dcTB5B#LAaW&44RRK3=L07S0ZHAP@/X2],T/,>>9>-d/99
4TNBG51:R/H=(DHPKVFRCX-X=FRA)Z75AN.</2gS[#-2.NR6VeWQPS@<I;A&QZG3
d.H=[]\OY6HDc<KP2\S)dc;d9DOMfH</_<ABYVL@)f2?)UIaS:JVN1Y-Gb4OMcHT
Q]THRZ:fV==0f1>Y2(F#?RQ8<,(YD.>,,P?O[7H&/?.RbSW]eVL[AN,E)+AR3bL=
=Z5LKJb__;TB69)^d:N4Q/;MQR<.gFg7AN7YbZ<^5JYC<,[(d,<g6419C+Q\Pb@I
2W6IdE-ee?_>O_]d(aPdYH-;X_?eR[UCc<)PSe(BRZ<.\P=L:/#,0G0K^8KS[Fg-
@NG.?#H.-F4KZ<=:UFOQZ9LD(JV)U>)9cP>^M:+K-7:JK,C:dX3Q(CNAI;#2L_P4
PU>3D=2(f4^;S2+-;FgN8L8=>B3_&G81J,(BQ#<SfQ0MSB47^?.gE;Xg2@TGeR5Y
aF[1;6V#Ufb_e+6D?7D2B\:EJ0NP#3+:V?@75\7,@S1-?R;H8JI6\.Z2?:::KWGb
cf_X.I6A+A?&K,7M3Pf?M]-8.41]I9X\R&Bc\aUA@G<f&+_M,EN,H1V2XW2Y\ERJ
9P2AeHD2cCR(P<KU:B\bEFFQD2MI<gU_eNW-dR8dTD=[<WWZA2RH2g:1]<gcIYO:
H5_d,?+?T.9-^aWEW,a(PgbQ6]W?)La=_BQV/IP9:M6g?X2(+7KgU2WR\=TH]T5I
aB?A\BA1=2.S=93PRFR\9]][VI+3.6[#@>)\KW_-=6b@SF\,aScSb,.D4<NW#^GA
_TN\UbNKQ>)Q,?GNMH2e1#):?\:D</;L1\3,fIB16Ld;-,;+TE.[NXE8=X+7WAKb
.<Pe=:1VQd@0=4b9)S@5<cATJB57RZN[R72HUK9X045&(K_GD147]2QD1^UgSc=A
/>,;]=gC96+&BF.W/3-U/S/^[/HGCX\:aFEQWU0OM]NNCRU1cG,+d/+^Kb^AN[g<
NGgF/d/b4,1,N\YQ4P+e2?(,?^JA<DZ;.b&#Sa/7e;REN<X4cD]W=83[F&.Q).a^
gP(#KU#SfBeRC)0eFM?#VMWBf2?PTfV6CZVJJ8c4SJ)-&?GOLH7<PQ0]2M=ZgF24
@bG)C6V5UYce>#M;E,<:CV6=14AJg8)f0T9c&fC#-#9L1f\05OBM@e1B@&W<Igcg
EeX&O(&=)R_#@N@VN<[;RSM\d9>W1N-C5O+;edHK-],HgZa,H)_(;YC\X;MBPHI,
bLW9eIW/dJ(@8a]fWHH^ZffS+^e-/3Dd2:2C<[Aa:T4+M@>XI6[:<E.gH;dcPW]9
[;aK;PC,XM6)CO/HZ#:;M9HOc:I@6)5fKBTKg(2WD,;(_;_A/+d&5MCKH[:#T49T
285cU@GcPLFF5D@g?0\K(bSdCF0<cc>:5)<:J#M;+e2WTK/&U/3@6OY?1):R<WLY
40TB5HbRML6Q^[L/4a(N#dQG731B72cT?G(@)&QF\A5QN&?+ETTX;GXJcQC(E&\.
U\UA?AMW69aH+XDYJD9.b7VXIJQ6?LDUX;(L/P75-7&cX(D)f3XR5N@F+99\b6C>
0HS2bEg;b64R^L11YNWA)OHL.:6K1KYHObb\UYF11EIHN.-bcVUZVRa?YLJ7bb])
:^a/R56Q[=OgRFV]PWH/2<M/&;YLOaMgKAR@]9=WYMO#.IT=O#KD+bGY3@)I6]2:
@LM\1CCd52ZH5c\A64V@_dD6&\O<LNLb9/PcdJN/@D]AGRGODDF1Q)Vb+VA5N_EV
D8dR(J(<?\7.JLS_M:HRFR3;7YBc/aFH+/8:\^51CPV94,7XQ/6Z]HJ1b<G2QTaV
fL;<LRdBR?ZW06\RG((M/O<;(.PfL@U3GN(58B>f;+\^6+d2QOO-WS]QEYK;HY,]
:gRVbff;+KN1bZV^DEIcD;+^W,62/SAW8WHP2X@KQ9D92b6^PP.BSF6;7)LRZaH;
>/3.Pd8?1/PC^SAK1LR^LAg4f&aE1@BO/J+LHbQAP4.7L8E3@bN0<K^2>9]E^]<g
eH<MbDYO4,Kf.C.gYed;aSTR)8<VZ@bb_Y+?XbA+J_>N1X+>\Y61W<gcVbOf73)F
01NaU<M4_4GMY@FJO=;#(e^02bLM&9Bc_)^V<C5^b,[30C;OMc/XP.]E9bL263b8
/^c1)2))f@S5.CD+]7NdJE@Fa;;MQ[WE5(e)T]1Q^9RP-E@_L;8EJIY-;=geY^4.
9.XS;d(7P0N[g[ARWFJH)W-Y(M4c()R.)g0125e4D,AgRfcE+NZP\Ja6/><LDVLT
Z6?QdE9U>K^3<O_5AT,YY6QW&15\_\3a/;WcRWf.2+W-5NaM96E7cR:/W+E8DSU^
OCM[.Z-[b]#3)]BAdCg?d]FIG5(^(D51IAXbZJ-@I>4(D?f:Q@dCdYUX[9/JY?7+
EH]0fPT0U8Tc0<B;H7V\NO4/2V7XfTB.E/5Ve<KV7=gZ6ET0^UXFKUC;edU70^M/
E45F<<5#7&gUMd[:EWWF\M_H=SNa_O;\V_#E._^c9/.KXQ]4[:\WRL:IY+X2#YR1
W8UIZL.<A20eQ@GRQ)[g?W?EbEc.U(T&BYVI),&:4AGGANMM\YN@)-Z@;\H)d01:
+9ac#J&d26O[4?40LPN/JWK:]\c2JR:MFBB>(?C/^TC<JE\]4dfC4XH\ZX:JN9-8
)E5-#]RggDYC)&fbI]QKNSdM;[R2CZJ&NFQ13+?#A5.3.3a,,K9E,g=GFV,XZDDJ
T)6+O81PZ:2Yd<C@[WGc1@8fV>Y^E>GZ^=AE&0]ES]7J6P+Oa2I6TaaG<09Q29RT
UJ76@>G5b7M(UL(?NX&^W>)8.Y;WUd)P,_?g8X7.H1RCdI\H>\Y3F-&CFX#e+E5:
#3_LJM17FMX[T779:[,V3;X,U=@C,)6WaHeFC8<\T<UH#XLC]fD5aM#GS:5bAJRC
XA>L;H\36@QV71gRU_2\aUBR?;G3@2Z<R:Dc)YUCe8g.>6,Me1STCg=2e3?/)dQ]
g8RB=@T.e#UF^-X==?#)J1?07dT:Y2YIdI@3[]GRLKHb\N/=c/\;DQ5Ib-;aX>/Y
0?df[;JLOeYD^=aPgQ7_0@A\8(f@QAcM]cdYMPPEKRd1M353ZQRM;eM5O+XGM-db
M6eYE-IK?5>:LVTUHVbXH5S-F?U[2f24SE/QTeL0,(fP>2(&.#NBfLBZa.b_(-cU
:<8dXQ,G&D(FFOMe;:KE&A0]:4C#Q0U\g82P/Z3^Q3OH@ZT^eV6IL:ccd4\38USf
>LP&&>V1?MK]79>YZHE-CN[N=BS9P[2SK))Sa:N?U+XN2/eF)[GMK9f/,_d.U#bG
@LBdZI.A4FRNd2[C1<\IX,#AaJ/(Gb_W/R_+<0a=SG3B8]C>[@X^c#Q7>EYC2aL#
6/5]IbPc.K>M(=V]/=Q\g6>Z1D^+UIBD9\JKSTL>8;N-Oa1JB>0_9.DeTA]+6aL8
3X-Bg0RcJ(AS[dJcAEM(gYR:]\:9)>5[V1J>/9OgA]2R9LCRQ^)7A&CWE>5e@bQ^
_64g5[#P-d+(39Fg,EVP>8<4d8RZTW1^JXJ/<(<MS+G9Re>P4K49=-)dP=e;9Z_9
9Jbb;)?DRd:^eV_E(>&-XSB++ga-@=UKMbR1HO</;+H.YSa&fb6ac<FUID>NS2-4
gdg8gJC>TO=]Rf=ZYSVaG,XYc4BWXA(BYcKcX3JP:+S&/X17<[a.85NW:=1L8J3>
)]7=S>f0dHQ5I0c?ZS+[HdYSS<QPZcNQe&Z(7()SV2?3I[VGG?3=e1:+e.8eFRMT
,L9\Pcf7+[#+b:7Q-EbBeLF:[T/CVK\1aE.Q,BY#gF9Ua>:[?KBXO>NF1FJ/ZBd&
C31&BL6ICPc<_dGfY2>G]4cWK:0B4&V7F@]HY+_PHL@3CG]T2[\SOF,>D>a_]M4I
A:dcA.b+IP6/^C36Z^-KFH7L?f\.T0XYJ_TKa-2&1)VbTU_D;-[0P]M>/9K+e_7/
4d;BVBQ2a]2L_P#,b92M^]S];[KBLIfbG^-#gbYCX,O+EFPZ8Q>Q.[LJ.&:^F_+9
T7-eU+e>>Y<]FcV5D3HO91<fdE-C^N=VGC0^<\LH+V2ga@2&L./<^ZFVLYd?)[EU
,X9H23cf=.Q,GJ1TYZH.JN_BHAJY>Q9b),<[/L]B)&#G\gf)G+8=.bd-5\PEMF6D
=__&YF<PCb:8U\]E[07,[7#HF<0IV:g)SSPKgX=BN6(:/AG@H]EG;Lb+F2:(1f_M
-,BA+JP_MW5f6gY.KE5c8W6+5+[3KB)^eAf2:,S(aWe7-3]J_9fa[G_B#Za1@[(Q
2PTgA/C>/[4F7HV6O[^d7TF^FVa(W=OJA0>G\2\Q;5D-N[XMJ72aWBKONYfT7]U2
2TMgTX-;A5=/]K<Mc;]KcP-1]M_b4<D?/e<Y:XR/#RHG=.ZY8?;N+bY(9Fa>,b67
J@&GC]a4OQ@f0OJ2d^8KPU+<1>7bf68J?Q,YJBW=Jg<2M=[LL5L/)^[M6CK,&fC,
GWP+1OV<>2(X;7Tg^0P]6YdeJgH+1+IG.C\[MN)L,BNZ?RKE#Y8P;#2&.#ZUYU;0
R0XLBAJ]V]aXN&:TOd6.(T.RF71384FZ]2>7=QB>U@;QH\d9ID>=\T\J.d3;F,GX
[-28M9\W4))babSY0<96b7#.EI(M,MO=.YD(Te=\.d[(]5f9EZHYBeP2J5c@=/BU
H.JNd4/H#A8Y+18@QN<0[/S]8I+>5TN#5b7S^+:IQcM1P>>Kd)JO:=&?#?d&V)1R
7\+LT148Rd]V,OL;ZF_#eK^7I_YJ=X,A_b0,B9U_/?N<?K^I;6SDgK\,H.2Y@-W?
Xc?E<]E01ZO:4D2Q#;>-&5.&J66ZW&a#]c1O98e?(E./ZR\@a.,0<HDD933>/6=N
M+3Z.0:aR?Rf:eSNYR/Rg#FP,>d<=90cfOO+(6TRLQZ(K_0bVMW\?cDbRIY3I7]6
=(;[5N7LDEe4MR/Z0LGE0QYB>cLIUcfLDf[I:E,XFV<CLP[T_P>S1bS+VPD1]V),
X6VE?UVSOZ3<3HDdc&Sea^8:a).>V,M6#bX+^)X1;5ZL(]967FD_#YVUI.c:]\WJ
[8[_A+S3P(FS/\:<@A>YV)(-_.fJ_SH2[O407eASR,7AcH44d<C]=JN55Qb_eK,W
C_XcJR1W2A6>V/)Ke13O;\Jf_XZSJ>NJ3Nf(8_]f(?C]-GSb.#>:T8^#UW?>=R]I
EG_DAGNZ36_R8(?4\e]UgS26N?K^4RTD^+O-QK.RbWaB(QE-G,;5A1BbC05IT7,I
4Y#N]XRF4XS?[XO,?96FVB+W=f&\=IXOIM;1F;)UWA&(6RBZ1O6U?AfF@;1CE39[
3]-<M,>Bc6JcB01=96b647PU)F-J@[cYG)2?.&@dA@d#/Ya2I2;D?Pcf3bPP[QC3
aGJ11.cJf.c8\L7EJH\E/AK?E5,3??H-D._g[#e\0HAg<=:DZ5G&Qe-OE&V]4bAK
:VAfcO#D(+LVVZ,WR;E75-dSUW7V9,30A/>@E-LRR;6dZSU/&>3SW)JeR_)dXQ##
TfF.MFf])EedY=d)CL.e--G#,237[QQ#1KVDJ_I.e:FgaP47,S-+N/;c/e+A&9,^
C0<Sc\A4Y6=1NPYCc_A=+dV=O9P2IF1f;CL.+:AIQ+&Q#R,F6NT7Hc3)gGMNONGN
9<.#a\&8?fTG-2MJ@V-O6;/=-MHf4::Z[acG&V-_<CCdJf-)M1;\ZbGAH-=0-dH\
4-R>,&BL>:720VfZ5egYdGWHY6_.0Z3ebe99/8MZ:L&FE5aH,;<QJ,@aQ(d6ebE8
N5JILMU^U+8&SQ>U/TW>ESEQ?YX5?]RIIF-b;7&?FVWUf(MFJF=3V<+2F,0U+8b3
;]Yf4X^XO^B>15D\PZ+,@OHBbFcL389UC4@]VeAA.7LB1=(#D2_9TAUO=(4+C[^D
^JbWS[QL5UBB(4OeT3cNHP:>\e:?=_I<F;1eCA[A.UZ&CH4HT:[]eJ]g=&)@ZMI-
.979-@(=U0>[bKEHfd#T.8\+bDC=(:=&9U[ANY&4Z8Zc+JTTG)=,LW(OAJHOc,02
V3>.51eHZKRWZ1AFE8#2J?&X8/VA1UE_G_Ee+(JPW9OLIee:6P8Jb3MS._8aOR^D
(#HB1b@@Q&Y&+f;UAB1=KD(81b2^aZ7EQd_O>JQ1L?Ca5&9RX>R_157/J#b^Te#O
5-(P0OL,)B6?DN&fWd4OUM[>)K--,g\U/N32Z8c=IIS<+Z/JF,>93CC:[IM?-,7V
+A6-4agFB;=G\A5W:)\Ng/J:g/_K.OC5aS1(M[QPdS.&b#@=F:^<<5C)fXI>W<=d
G8J0AFK/CCTZbW?cEP.[=Z8;bAg]\AFJS]8.GeR55Hb^_fN<b@4RFPQIH]]2AFK(
MPI=],HSC\)AKdZFRB.?8]@:QPK[d,EF7c2\0RXFEQQH5Q15O,(b_L3I+NCR-66(
0_=;44aDCYCG317UZZWE6-O,?A.MF6>FD:R.,ae4(6Ed)ZO?5b]D.cf])XRNIL9b
6Z#4;7MPX:f-52;=-6,]C9LR78T=9.=HLRV9UHQFYX4ZgGdM2P=R(/_ATJc;OOe?
5DMb[>OOVFEG\9LGYd+bH&B2c(HU>LeX2R3TT4MGB<ZDZ;/8;8=CU4^3LO^>V5NJ
#+VW6bf\e-C-BCUKT/6c_/Q^_Ga9R3E0/<^GJN2=KBXA+PdVg1N6QHLd)Q=>(bO6
PS2SIXK(2TT+I^BbGIUX-^-]LA?Q4^#U1dAISfZM(GN:YU+?B.BDaF4+D<MS7Df9
[5@\Q>X8[<27(\-D2E)(7?_:/LZ2^8,B9I@T8E#QJ0fJUcYgY]64fJS,9R7R1PLf
F:E61K6=;4L[UHCL[3=9-#E8SW,8YLA_0eR9(/:TV>FQM_AMH(5@dS;C>H6VEOQH
(@gCfEW?YHG0UObA=(ID[B5&RQ5cB3]LW;UFag71[\>ZR^JSL1/)S,N+<b&:Z9&K
<?>]M]4+=:UWY/f4V.XS,)fR5:V[ageD)[T[>A2WcN<HAM0:/:bf0-XE(4fZ-IHa
UFHHg5\dF5_BfF,X(HE/gAFU;6_5WZdK>HFW>/^Xa^dM:+/N91Q2fRM<b:?Y066#
U[QW4[;@#,gD8.d>,\a\^W_#)2X-HTc.K-XA(H:&&1Ic-R+M=f^?C10Q[)+dbV>=
;VZ5gQ5<,DOZZ/HBbLHfD_eJ\(6g@RZYePc6#)3dT8:-F/bR\_]IPVR0b-+#d8ZW
E[b8dOd],D:Kc&9?-Y<-X#=BGZU=N@N(3Ig08JX#HYEbMa[M>dZBUY;GWJWS4g4W
_QUBUP[G,=)ZF^BT/WI([SNHVMN(f+@<C.EI1@Ka6]?8\>.:QWI?G]7L<0>9d.?c
U;ge=G05^01d./4Bf0g+d?+HL=RJLg)8B[;_WA^?GCQQ[7(C@3.HE?V4&/765/;B
@g8V4G2AS5JOI?2^/HZUWSF:1]B2B_Gb//LHN(0_(4ILK[GYMA@.2-d#Ib0eXAI.
#SPZB?MVG?]D0HR]\0\&N^M0#.eaN-E\E&BDS2b.OP]QCMG.7?]1dY-=B@^J=1&5
+9W-<(^YC/<OPTXQ>]DOE>+I)ZAg@SdNSJ_M?^E;\Da[6J22[H\F4^//-I@3O2g=
D4^B>UMJG_680d6[K-,V4BQU4:N1YKCR,@c_&aX:E55GPMf4eZ7RBB60[Q&<7M0;
f^18SO^E[FGE7:L3V+bMN1S4&OcKf4^1TC6HGg4?VE2AJ\GLNLI5Q)5X3P=+fd3[
7.TCgZK@dDda\3>9Ib+-eT:855RAY+Je:]@OOVJ:YMB:S<Q,(<>L6D]5H>Q#H)?H
@H2cVLTfUY8)5P8>RK\M2JI68[M:gJ0K-ALf=M4@]ZCGODOV:[+1M5dQC<]ZF#cc
UAf5/+g#LJ@cD\HKK&<[Ye&J)),_P6TbBLRTWJR+C0>RC@=CV35c;YLbD[;a=.8G
&9SF0/TaO&YBGRA-4FfAHMZ>7e[^d]E@QSgS:OYNZ^958\RN9S,DT/@6TRB=R[K\
g5)JDC1R[?[3QZCGZ/06^3Vb:R],J)a5-Xa?-/_JL(+]7)8J8&)A)HF)SOWI(@&3
C](W_AV:JUG+M/O,;K/)eBDd0,48&-KUZ?1bQW;U)DDK+>=PUdTI0S]Ke:a2EK6C
&]B@TT_9Ya]F5eJCL9bfR(L6DTbbX&<F<I+2a[WZ.[BK:S0,,C7KaSKUe4]B/?#d
UC@AV.Y-)H6&Fb2e+)>.OZ?Pdd6OB>KUG9b.5&5/^H^J?IJ]X))L=g\O<#+,+g9,
8YOJK/[a=>\Ae4FQ@:YA)IQbDCHeP+2L=?f:GfGR=_;K.Y7P>IX(Q-6Yc>1dV=@8
.9(Qa=CggPVCU@ZgAc3=f&(Z(I6>U:CG9W;>^5/5)aNYS4S_/<Z^@_3>gcYS-\+b
5LOMNYUARL8+Z,B)9fM>-I5dD\G.C>C<(G\:(Ra,BF8GeaH9aB;6f=\H8LH./1gA
e7f+TG/KR?fDTDGPIf_B>5#cMOCXT^04QW4OP53I_4S,fSKcVP#(fTUDODaL/DAX
O-D.Ke[O,]G&@a:>gVc_E+GW6I,B;7_84W2]ZHST<W(R\=EfR1bQC1)U?[WcE8I/
=g#g^,JL?IOL-EG,V5ER)PDJ?D@M<(GBF]XBMROGF:^15PKMJ(A^Ab@aU\E\4SB8
+agGT?GIPAN9LMBXEe&4^/+]2&MO=\^>6;GCD8RX]+dTBcXZcY3OC+Y5\BLFI\(-
P;?b:U,Ff<.)]B-#.,V0fPZ3DTbM?@FTa\_HTeGB[Q9P<J2/,EO\5RbSZ15gcWVJ
bD5E:NTHR00\0N=C@3_,I.#(47:TT_7I6Pb<-IJF^Q<P)D-NR/U.E@f/?8>?]\M0
#8PZc<,6TWWFKg93LNP+E85dTM&?(,aP&b@^N+1#WJFG?,89A6->HZ)=R3#PX]da
F#6TO[cB.,J51_SJB?,;/A>+#B=[aY_FL(WCDQENPS@9R/[.BfNK<KXRAeQAF3ef
I(gXGe92Y=G31d3=R).6ICC+9Y8.6L<0bVRXe:L^1bOFP-HZ?90;]U<Jb9#L+G6A
OL.O0fS#=c\\ANCB7;FgI_)F1(BLKQI\2R>,HLd;P3?2^bJ68\g_[R]d1c2X515#
\/SeH5d,KVUR1Q3bSUIV@LX@8e9\06dY?\&a&\2\.a8(H+8LT4#7(Q7@Mb3@B;G<
@O]PJQd]=-aO\8aE(Dd0CP?VRFH2gC)SRg97E\(/>GJ\JOJIbY?4G\V+.eEC:IQ3
E;AcEgXdDf,\NQ9Y&NYc&5^<VNU\>dCLcSGAc\ZJ+>]fX@H_BI7CfU6fdQL,CM/A
Qb+@(9=f@P^4C3B/1_R1(4U9]KV;R4M5.5dLaCS)]>27=/eZ8?KAG=G6(fLRF<cb
.S[X>UFVe.UM\IG0;T^(.cG>/OAaRf:.7;)0_+LWJW#=5LE/#L/[5?HT#;CPNSb)
(NXO4IcE9YgDA?(CU[3MNX[M&7K&gb8BOI,E31:<&7_d0,#BKPR9fNf6ZD#7/[3;
f]09eVb;fH>?gb8#+[_Td8)91g@60REQD2C\^+2:(8(<^+&<eV(Dbd@REW5F+3Ve
Z(#IE_LAfU1_,OW,];&c:XL(9>Ea:;H-P,8#LcO4FdFfZC9N6X0)A2Q;:VZVb>A0
,Cf)(a,?7Jd6:DbFXJ7[\,7EIU5EDc02X0DK(QCBT=\/_;=/DZ94[_QWGa7SDUb]
[F(31CeP\+P[:&B.0JV^>-XDU47[DfJ3@c-Y<]=LCgAaY>@YCT(A6HJ_4,&:@(9P
FI#NN,;\B]a,B@B(LPTcJUgEbKgI>2RS^<FMVK7eH8OMa-A3R[&:V/&&g4dHAB3I
J\;.X.H>NT=\]-&\HIdAb#3XX5N9/+WFD?TU/=CCFKON\1dBJ9C-d&f(LXTfM_C)
MD.W8W;15H[8I=\e.SQ(ZEWe<KUPM79]T(d3>.B-5X-cf&C_PJd#M66RJM@Qg<\J
[0K(D5](R#+a+1#UN_V>21VI+:8)D74-#;@aF1Lg/O2(Tg2M@VK>/8\N[cEM&WYS
PaQFA[EZ(A)-8ec>+B0,S>=EPJ)&L+/EJY&:P3#6;c/.a2YD[=;)XO]b_QDWHd\8
SE:6Q+X:TWEJd33e]e4;Y#eHA26fZ9ULC\+U>N[GB^O/,-P4<J>#A9c77^M#EL[b
[,dS/0M9^PX3[<.8Ld2c/81:dcQZY6BdV9BFA3B007?+T,c3Z,\VR3bD#Pe-4gUJ
)cb;CRFP_G9WRCP-BPdP6d9&]S>](Y3?QNMgd4Q2YB;_YE:SMK&;G)>CcM#,+6KC
=6#/J>g(63fab)(KI[C6+V>ZRHFV-3\AH0Xe2K?4H=0OHH]cH=M;+M=gAf_]]E>U
9=Z_EK<B+Ba<-_f6)7Z2BdLFL)bXIV5>WQ6/Uaf]DK2F@I&8WUTNT1aVJHe(\d]3
WS(2Kaf[LEMbf(NK3fa_O4g4,S=B>cFF7-Q#AcT91S=b=1MY8RXLG,?4EVB9:<d1
R]E36U#<<(A(Q=5)NXYeV?[cVEJJEa]fGMe-7efJ_\L5I]JGA83a5d_8M[S@\)7A
&N=^-[A6M0,_Bf+JcX=,8-]QgLB.a9JV?@acNa4g4W7WN+1dSeX3U^;,57NA6)-Q
,U-6&_Sb(;M=@HT8O-b&V..\Va&^\6PF25QfA5Wc2<Z;2#5V]23<La0b>-/TO[_=
0F+YNQWa7I)7R5X1:^L:<]0D&9E94aa6HDL(E[#,FI<b>RE8\d^YB[#d-QP(SQMO
=Z.3e5b;VJWWfHV5X\[NTSc(MO;I=S:1bX)1K^eD/.^K/WR+J91UcbCa/BO,[N2g
=NE87\V;H_/(Q@gg+_UGQ([SX-&]f56H12KE,7^C(Lc#@gKDY010C/2cRY,8M-3F
K/<ORG2_@=0Cf0[B^P1AB<PZZ2Z,a;KR)?b#@F/7^-\&cf54KO_fX8Raf;M[#I\5
A4F=5\UNQ8e1-5TW\.XQ\OS^AgN?RI0O&L^P12[^8#8[BFFU--dCU?7S25.E-JdB
(^CX?.BMCN,BMRO-4@:ScG:ScUCYUI/H?BfggD32b?CG6.)0\bX3V@GH1.I5\LB@
)NU;G:E@;#9>7YJ[,);CG03E=WB+?PM2>[_&RFA&.J2J?]25Y,g2TOK&ceM^K.<H
R3cZJ]<SG8<5:@UEL;3]CGX<cf<cWDX\1.\#e5<<0F?0M10WB5<E=,-ABGbf\4J)
g9^12W_<K6_8^.=H=/@AXaSdf4>KW/bPUX/+dgEJ=0_=XWEZ_JSY,FYUDG5LZJ3P
C[8LKIBKfB0,3Q;PABL#?I7:H;WLER<b8gb,KOFa16F7>3OPF?ORY5bfMQ>7DOgb
R4I9L^SCKXE5[cM>B]PS\?5ZF5;A<5F5Z92B(b@5L;3+\M;^^IT(4)P\\dP=#XYJ
_2:_<KH_ac=07P+A3gVaJQY-Ffg?KVObM>DfOQU>d=Y4[W#H>T+_F,?6INZCRTJ]
_#C/#^aBE7EKbF(&?a</U=a,SJE(N8C-M?eXX+]39M4YWMRgX?\UF8/ZTNJ^N06C
/0EQ810:-UR)8;+PY(>d@>;3M#>YX50LHE/-&#2,dX6U_PH:C:6ZL>]Y:GPDD?@B
T<3c63JfX]?6AUWTa=U1a</dB<_DH0bIJ4#GYdQ&P/J5<=Q\V\M]IPGTI19TNTf0
49M25J(15f69WW(a:aEOL,4]Kd+\=9G;N.7Wb/eN3UUUV-[NSUI8LJefM/&M;;I.
5c[NI,G[X&8K;S=M8[B.,a&<^-=+Q;]EUBB\gHIB\MBVbFb&]CC/>G7_)&N&_QNC
@?4T/c9UC+Q]eH4.^8Ve,(+H,G][\#QQ]+E^QT\RSSF.::bLL4OTSfP)4F0cG^9P
IcRSN/7&fTc-<&]DM@,?G[)1@&R;GG<UcQ&MWB_[>^G@6e<,N1Z/40.&A](93[D(
A:9Q;eCJ]NX#U?I-&g[C<18gA+e=c0Kc(:X4Y#_dDS+B[_YY:9_L8>#EFG+B(RD,
#>a]5H&]N[_>L5Y/Y#Lf4XS>.-Qa7=5F_edO&Kf.>1,1DZML\^(e,K6DZ-Y#;&6[
eI49U-S4,#c>9&[6]X=]@LAM-:+]G8>Ke(7S#NWNF=TZbH[ZU3J]X2PI=KA(+Tca
#H&Oe[8-?A11U-V1XN+_D+4D;_G1WHUU4Y<>[d@#0:)5J4H^1c=HIVK)((+B=Ta2
J0),J99Xba4EKGfH/1SWW4F_I7;M-8<ZBIT<U7Ta@V^0Uff3aL+f2#Q8Z/59ZOCU
H]L_bNc0BZ5C&@BX8A76>0C\R<XJ+GHVO0:UX(9B>N\eXd.cFR9\:=2:aW/-bgV0
G(&B6e&]7\3QEPI9I#D4#eM_I[+-6G(d#.;cNTVK0;3]0EFf.D>8e.<>Acc8aMP+
c:FIGP3]TQ@&D6eR1DE-P301@MAL:I1N0(a80DF>:9(b2(#&.IXYAV9I5\M]I/>M
e<EA0A8;.d+]X3(cc1>a[,f+9_Hb+2T840a]CMGNJSANJF5)#@TW3VX\Af2LKMd2
GHF0Y-YAAR@[0CEVKOF=fDBSW)c[)@<LO2,MQES0PD0=U_N08YFTfOX4fMG_4V:J
I#dcD3VLJEFg<Q#<HVQ#9.?.adD?+Yg6HI8<O4WcgGaW15[)T;G]aec3:(2c>,7H
9,M(EJK[VRKFZ)E\0669dIg\I]O8SfK.UX8\=1(XYXgB2ETUb,d)c^Dg3g??(B@N
;&adTCbJcg&fB^2b3,(0O(fCa1+XE/T;#/RebK_fXcW)MeOUeMB7.T\HMAMgKGXH
A8^JEb=d.+JV@NP(QRI<+V_:_YNG/Y@BbUH6f/S+)IC4Y?d.G9McHdL6FHR(S/]U
4&T63Jf^NQcR^8JC6;Y5GISBN5F.\cNQe1cU)EURY7?ZJg52TM<TYg\9MQLH3=J<
ObD?YJF<<.EcUE-8f]?#1DV9AaRdJDE,X69_6NU#b80Ub85NbYU62=(5BK1fd0Dg
Y(LR8KeJ;cO&]XU+[\N27G]/1gLH&E5SY-I5:]E2I^6WV,S1,XcHUDZcZ&6Se=Eb
W.g?c0>8T?+(_ALW^VaKXfcL>P_UYH2PLd80N(11=e^g5I.fA_K//<->/BNME(-U
K-5>F5gLA(?R+9]Q-U)>;I))<VBOT8(BSKT#4N4b-#<@NQ/UNSI,VTRgEba@HJ;K
Y(-DDS9S2&.e<bcJ(@M\@@3_YDLc2ASa8T5I]OV=_?.&R]EFTT-KY/=G9N@a]gP7
H9=>[(]0,?]#LW#W04??87Y,dJ=UWSMT(N-Y27bQ)+JfOH-MX-V.EQN\VT;N;LS^
SH?Id).<Z7.c6?Pf/R,#Rg.c7M;KWX=Q1SD3d0bZ6,d>HSX[79TL1e0;L_4Q@^;a
AGD9B0TcQN.J\T)8?g;L)]><EE?AE.WOT(RGb@C1Cbe^;b/]CV(1,(HSOC3e3,MU
5?W.XC2HgDPBD^XLJP.A_O\D-HM9,61G.a-4H7bZ@:R7LcCT5;^bNB:4KE)/M@9]
1+90XC=X#Ic>c&^_E;G\/cB^RP[Pf8,-0>H9NQb6[]e4XN3Wc@IGV]NTd=H#K]VZ
M20=0N[9g5eVA[YGKS)6LWFe[f.9R^.8fLY21]21K0(Z03f3[51CG_C630+>PWNQ
c2f9d=QH;&D3+dIc2dJ7bX2c/GT/g6QF3:L47O]\EW0dZ39d\Db,/2RXdV7:)Z>c
P(75eVRH_dTfHBX^U4-WWLf1;a]Pa=O-(#98D-G#,?Wg=6TEQ<R_KT;)K4fLJOE<
LbL=PgSgDH(QdQF[cW^FNI5,MG46C(OaTC@aJ>cFNb#VAI6)@AP_)ZRY[=N0b:Za
KNKD;:)4>dE^bbZ7SBZ,F41P_<2&OecN3=R^LR6PSK1XYX]#@f-2X??@_DOG7\7C
1gCQ;c@ZPB-/IgR3Q3]c)&aZQDDg;+AeU1:fMT?4&R:BUP5H/LN@g@@,J5gT6[CE
75WCW&X5)=)G[G;]+:TTGA/]:2DN\ZHH91SNU]S?Ye8BBd#Y(GRVg;M3&:88+RLc
[=K#,H0NPZ9FE>I.\.FG?YU,82=+#JUKPRG^T6aNB;JKdM?YN2:,J--VD)3+Lgc9
4#OD9;_-1a_8ZGS:MRS<IBRM7/Ga;+CXP.Q3FMY:BQIaDbHb:1S,DFMZ1.T^[KXg
94A(0K43FNB>bE-R296YbL#NO76&3SV)\/,15GK.SQB0R;:=7HJQ),AIcP[H^7gb
T6fUTJ0EG1GWGPgX(@CO/JgMKCJ>3-DR2eZB0?dD99EDS.>C\&[\X;,1Da<,YQEZ
_]FB+B.2f)cI^\XE?(8MS:]C.B(\SbG6]g^fM960PK-J(B=Nc;[aJLHH^?5.VJ@G
I_F\cY=CFR\IQ.FCVEB6E[8^^_aD3_\-ZM(/+0@[dbO,5VK8M&DSRcB=CO]HKYW^
QZ+g0Y3g-\b8EcTC<BZQ5BE:)U++G.61ffeT\W,,g?JXe62Z:O><YO(;BfO<M?He
#-OOE9B1gf9P,OYHOPQ@O:/CRMR+[Za#?c54\KZ)TQaUgDS+FM\V0aVG#_ae1b@f
BY#:Ld.b?/Z^_aPMe(OWEH4(U5PBeJ\L:[KfI;9eOMCE77GRe)9GFb<K=1I/]V#]
RcN?[4FX\aE1=B9=@eJ0GKT1@+.Z/7.-B1cT@ZCLSg9[6?O[6dLeBB5UB/@JALU>
FfgL8cJf_AO&4:M@57MRK+HK+0C-I^A/RG;PK9RY8?V29H<ISJ1^@^a_WT4N6LT#
9QX?/>^6-6749ERUS:7Kd0WR1)Y4=OPce/cZ8:0H233@;(FbTKMN4Fc_R[;?9Q6D
]D1X7>QSKY<d\-eC.g)B-I?dDHW)eNIZGTK.NH&CRcTVQ<5KW_I(a2:JHb>dA^1G
/fCJ9[W4X(0O,&c57H)7]Y68eRM=g.6]\/CZWLNMVW#M#_E/#NE80]=P@_bQDc,;
JDd(M/@RB]3UO0FQJ\TVJPCIO7gLW7B;a^:VeB+c+AB3#KGZTf=EOBZHFARI6NT\
:caW=5+B3b:K-]V-XVHX6Mg\O+aBRdWDQFB+^KS4NeQ6S7=]&=65[c+GQ=0[>_X.
T=+]eWP\3A\CLYfa?VOegTE3S6T5P)\O^BY1_6U+G(0\.0:20C,C>\IGZYRDJ&WT
aGJ-?:GBE\F]1g?Z3J^@B;fC=#<T[_H#94F96&80b/c<K#4QR2.+/6RL46?9,D[_
JV110PY>)3YP0ZO+^R&6=b-4__\[\:Rf[Z9gZRL(X_J9@3aQ^2;;dR7Lc=M<J.=/
5GE5GC4c?A71_3Y(UP_a685XTH+],J)6cfJJUTUVVB_DI@>cA[a9WVTD\+?:CZ^Q
3)[;fF]@JIS&@1(SdUY1ZKR]7c-9N(F3G2]3M]I-DI=XK==XM)gOQVC(b^F+\^&L
#b,5)V+J5H&F(C<VR<##Y6Ed+21&FeR_)dTD(W8;U:Xe-JR]L]ZULeX,01eMTSdY
fM3dAI#O6:.UaCD(E4V8CVN:>I^eY(aU#a.1&5^d8;0L=5cP+OA#8>eU)PUP;89(
R#<6(R_43HM?=[@)L-;>2#?2KGcca?H42KdVd;5<_59G.QE1(&HaC6L-=1NHa?S3
>E--+GgTb2>b@a708FC6bHBI(5\/J]?J3N[eAP1:M((dG<G;@f;N>F;W_0UH5\S6
?D?=^9B52#DCC.JJb,[>/(7SCe)^@M;3H9KJdM;22dT2O86TF,Y8Fbf\4fZ4NRL\
T?1R^<(/5f2EB#03aNEe@W7;f-U=[<gT&\;>(?#:cc8V-DVN;61a^+/c^dGI-_S.
+]fbGHE.]=\BJ>=gP-)Y-D4I4^;;\4?d8>7#9EEO2^DZF:F8=\A,?Fg/\8aTCPU@
1<//K3g5I9=FcU+<<feEYKE49#H88?5L.dN0.YNHdP_CP=-3eBZQeQ.9eCH+bNH^
@,aKCPZPdHXf:cZ)6M6_dD](53OR:MEJF(4.?@:I(ec#G_c^_N92]\>;FZ-7;IZ-
aV;+^HBILR5V,S7LA86)7)I[0bO4Rg?K\C]BNUQcCP2#6/1MM:Z3UbL+HY;20UGR
[VZgFfb+E;/S+6<X(+AIbJP4G3RXG=]d_NR.;2ADg\BbJQ;,;2;T0X]F(fI0#Z+6
#EWKMUY8\c,<#5;0P:7@\MO/M)J4Kc_8W95W/46_118?\6B:P;gf;9Q1>dB_;[E@
DW\,=<T[g7[Y6HS[E#9KdI[8A659AQ@bF9Q-#<2OTM:M<;b+[T7O:b_QP:84YIRa
++eRZ2([P=;Pb0)6G.W5c=7?3XR3-Q^WXQ\eLI^:2<FN4gfM;?&[8Nbf;<T1Zc<g
L47?O=&7QcFcY8W]ZC;02OG,AO,2;I/.-HG_5ObC-E?_>[_P\4:,Q4Z8)H@<D^_5
1^Zd=[WReF^FC2^CdC\7^>YC9B[A6ETA<EJP,T\0U?T)D?^@BgMLIZ1&f156&N@Q
eR6[ZN)6T,Y[4P?R:eLg^4(GC1YAM:<V\BJH]BgG&e^;Y71VZOCgDD-G[J9Yg0#P
2ID87=68MdXASd9aRH>2.+TeUF#Ea]82Aa5M4L-I-bCB-Jd6)9>,^C9VdX^=4MYD
HJb=PI>4a&?UdO(cE(;(>3[IRUTJP#+,&?IGS]&@2AOSaIQ[J:>59^(<g#HdY)2[
=MYM.FKCU61RQL.R@EeQH\b^g\>8AP19I::W0V7?]OA>b@_<N_5bRB8G>#Bf?\@c
^ZM@N2[]O/fP^2:QVb/X\F45&/E:-/GC6<]B8>dB]=Ra\LNgUDHb#A\)814EX(@[
G[;81f&A>+<]K4CC5aE_\Hb.=ee\8+0a=YPVFHW;Vf36R7ZOg9WL(\UKTf1/gDId
XIg8Ee&UaI[/EUMaS1U^[/Y)X/AK(I?G8FefMXS-c2>9B9PLKe=11Dg@YO@gVe(:
K-FPH@gJ->P0#3O7Y]Z]^a949.)Y8^=D(EI(^^QaJ2/fQDEI9>.e-NdB9e.OJ>VE
;.G^>07eXKMS_ICNO[29gJPcf2B@0J9Q/b.;IGY>9<#CCPaIZaIID>Z,7?4_I4O<
beV@.FS9&c_U[=#RQ7W7I>8>HJb_?d&&DdgWA,[=[37b>aG9bPR\WM+0@a&#L80E
A3))>>OH7Y3c)2U6W^_dI-.IB<;SSCT(VPP0YK7/K<L<[,<bQdP(A(6&c0Q(\A9,
7SI,b&<3:D9L>;X,V#e/8S=;D+TfWg\-.Pa&d26DbR_,c)LS&bU>=VAa7Nd.HA+P
dG98&7#\3Z0E.2FJQNa?.Ab.G63@f[<aC<IM74M&77^:f(SU>c@^:-59>Ag,A+1W
DU=T--_?cZA?P?2Sa7B[bA+FH4V^e#L8d#Ic:bL]V[EcgVcfYH7;gdAOC<WR7YY7
HX(#e>:L2LV.Y/O=M?IZGI[IG(W_W=de>aebbI,d?C-,3PWOG0<33-cB93J1W=V#
<.\:fddN1QgMBU9#+J2dDTA;._C^CIbM_JIW3Z/;IZ(dZOgATUO&^:?F?Z2EE5P>
&gaIcI;Z4MO>+PZUDI@ZMDT@;.D=/&3D>\gQbQ=I=8/d#f<bB7VBW+Y>1QAcVe<S
U4a\<I@[C3VOITXKYgP^<JW73BLV>e&7G?;J2dPTLD\c\]b3S,_1ZM,=<)A/16YI
1=481_4EKYN+0RIB__X.8:?PA6Bf_VLe&??I2)Me&=.341O75Iac1Ea&ZGS;WV)E
3>ZBFVBHX:=]8^GK(7VFDPU0-\[d<U,QYTNL+Ad#GV;Eb>NSZAe]HJWI(d3]#QRK
#g6/IfSfVM9+W1(9K.E.>I_EN<([_DeCM7VR&+L7B=A.O8FT(F/aCX?HPU2W^N3#
6:FFQg=d23d8/gdP(Z_/3ONC=2PM]204\eY93;J5:B8GB&;C2>E[/2<#gb_cSU01
P(gPKT1),_Kd[,_&J\bGLW5#-d7VI0[O8QZDQ2O[GgVA9W[:7Raa2(1STbZ[a/Zb
dc@&0G2cW2QC_F>ZW>0e9_AWGS/eEb83I?8bJ)-(#5J3B.IH6.<c<B,3.#X(J8?#
(]JTHW3RF=9\;>J^6L+QAD+XWC9E&6Y8YX1\2JVZ(,d:cYK1aQH<d=;gf[/POYVP
U.b=g=ZKfX3H.GE3bUPG[R9Z+V0M4N6NKeCYP^>(fJY9+:4e07<&)UU&ZL2a^-DC
gB..2,M/)5GJ(,1SU#OP)gdIOQHQfZdbaV=CRH\16KD:X<L)>f45WEJdZa>7D0=a
0@8bMO50MJAZMXIAQ&M-5<P<eSOOF9M^XIK\<8)#d2fbU(#?;;aM1\=g0&L3d4gZ
?f0;2/gS?,T?@1bUaF4=c.YF/AETXE?eK^O8H82\MM7&D]0FI]S-WW(Q8@T;0>AH
J26N42IaU)I5/AQ1@gODJ:[Q:g,P-FZ:.PX/VbCWS^d&/8<J@)Gf_UF(,7S2^:cT
Y+48cK57CM_/1V\V/,\YV)6OEd)7PNT78H)93]^50UL4-DQ@\J>9P)]NA3-c0.^#
3:=Gc,;YKe@QZM8d@+&HW6FGA0,&WU=&JHW8F]aFQ6S&>\c86OgV?JQ_Ba]WESU:
\]b@(FE3^.[dW9477g#4\G1]6.R@_,+,2@F:N\HgPCg_9#EV(E=UcAB;V\J7#0Ob
>DTEa))fCgX@,ET>R5gW(S8(\3WCJ/3XD1?FUU#/X>:1:FL.M)H.ZU=R:/8f[4F.
5])8N\E;+I_7J4C58PQ5QdT-;HK=)9T5eEVE+Ra8NIIT2.Ra#\H#^6fa:MA\=FR4
#=6gUZ85K7>X1C&]MNTM+SJ&&25S2,[,Gd78O,=SDWW)d5[A-C(.5C(,=.468)HV
OA,_)YfdF+&(98UL[EZLcF[80GV<0)g=<3\bBQ9#2g3RG)1.H4OQO>gZ.N+,6GG:
G27P:EaYbf0A70JP9G04N_ILO.]1=gd^gB&ZQ@5]+EgK[F5/L0QIIeQa@bP+_^EG
JIVWY1D=[E@O3NDa=81J@6O03J+gSA9/YL0/O8M+F\DPP^<CC]C.A,NI95c&)c:#
ALA6F6\8e]ZK[J8HDR^=bH.8@aG1&0,,:31P<)(]cCJ-\1X1;/;d-:S&\\=U+VbE
EW:eJY>ffP[OV9^:VWW+N8b?H0dU>WV-DdCLJ>[JKH2?d8R)W<72VNXBK09f;A-=
[8##8NHD.-cJ30<;4+K(2c(U-;-VP1T@e:f;[.03F(>@36O6G_fEB##?ba\AMgdf
KFcVdWDS6^,]N+<#A3N?W^BH)B+\eJF:;2)CAUa#8Vc<e4L<9P\[[GM5gSEeA(PT
S#F@AEaDUC]gZNO]78,HTM)f7HIe=\?<&(_PEAbS.\:b2/KVC16]@VcGS5fK8&9>
[JPR/M;f2RBg^Y3D=,,YG1@,4Y2UI(@Se@,2<?#/@RV\[]^G8W=U)^4(ZU]fHff(
fb]@_;]]Hg(#(@];)VRGTP#.K^,CXRM5A^<3:QZA/1&:P&O#N0_^PN3+^3296#D0
?E&V5c>VLd7EH[WK8f+VB<?dd&b&OEWG.FZ>16A>2LFgU5[0)P9;F/4/H;#-_6@F
L(9@DO1]39R_XdA&[A+UDgdX+3_4TTLFPH1DSP5;CbLE7-AF68,XJR\Xe][J3=/D
[QA/>2ZIH#>A4?:Z[YE]:d&Re-D4>H=^Y6[E@K3_8-#]V[L2M.3R\VFX5bTZ0MUT
.Me;.(<4?1fIZ9JO=8]f<,8^)Ac-gcbGa+1L4@NOFa>S6=f]S-gNBNR4U+/5[8b_
A48.3XTF[CQ,JEWB?HM54Kg9\28WR.PLM=fZY?KVMb&UBZ3I2]2HQ0OI.;,V+5OY
g@UKecZ\L1S@fM)D,K5G4.SK]#?\@[.G5XLN+O4[6M,c4S0[](/SLHA)VJDUWb7=
fY_SI=fJDcN^B?#I/IZ0YSD0=5HgC,WRg;70D8H@;PDNVI8geN_6^(#,d_<]O;Ub
b0=N;FD8LELA>Ue(L^7T.P[C2?\:<N^JJDaaf.]7fHE5)=76A@c>?[XT-]0^ES+]
Fe=_bUa.XbT_IW>5QSNb9O(#>bE_LP/(4&S1/<YC;UI=)IaQ5G/M,_._J+<OV09S
TS_,W;JCII\8R&A/:Oe-)d[NNOX099KU;]0S=369aL8UQe6Mce_2]MTR./3Xg1#L
RO55JU--0H952Z]6S22KeZJcZ@=\]^,2T8HU>U/Y=V924@WJP7[@3AMc2/\U]47e
A]6\+4>X_65T(U/dB5H^\JK#&\Zg+bOO2NedEf=d5g]P7S<G[9F+JS>YLdS]-bI&
-H4_Qf)\^fYEfK>F/^Be7@fE\5Y4BOcIS(KZNgAZ-LB5BVbRPI.e>YJ<_=MUACRB
c+]/56OgDgcDa1G94<7bfCMF>B_?cT;9?CI<\(OL\K57]6g><D14OSL24]G35f9)
TH(f:S0G@7L#1I.Q-?/Z<Z\@9_+4KD.Y51T13(O3WWaD@@YTB.]--PHgQcF7YPg-
60)2+e/UQ<6]VZ-6eDJ^ac0WLYdHX6LU\f-(SYECU823+:Me,JWV^Ic^OGgX(R8@
_>EGC>HV9LDZ3+77WHL<T>ffVB#E5<B&#,JNB5HK(A.P\LQP(E#&MBXL@8KAH+0g
&1Rg\#K&NV2Y2AJe,LN54@OKW(24aW@>_]JVDD-R&W@Z5B?/_\/G>bG/9T>BVdXb
RW>7,O(OG8,6N#/S0?U__BNL18DMcS+/a>Df?T+BYC+5SVO6+dQ9EQBG<<\^-]&c
b?fd6WW5L860F\HT/c/J0\dcBI?H:aPM@ZG4228<1KJS]Q&=bf,MR?&gSO=f[WAR
\aP.CR3,=3S<7\FOVZ@04KU&AB4PEX-E&X;).TW=^-D:\(+f7ROX2e+e4(0:PE&,
XP(QZd3D/7N:acf\?MQ<<W[Q,P,9-HQ5CK^\N2Xd0g15gXZ?IA8#1C@I=BMN]X=2
<9#/O\7Y]?aVU[O7DZdIG24[aF].;^2BY+)<#6+#]K3=6&X;W])JEOSA)PG()Z#.
AEE8=W<>+V360X):;QR;GXL7W4\fPFS,d.@Wb)3L6);+X67[_=fAYLR/VIb<3d3W
B.(?cR20LD-b^IE4a68.J/R45]^,9c4Q@B5#;K8)/<NK_WH=a=WG0UYe+.#?(QUF
X/HH5e0HM5?U[68Q\3c7S#A,M@?d0OI^dG^_^WD1dR(8X7&A6B\_[BT+Y0I:R_3#
U87I/:LQRFb>\82(C>P7@FcZ=_H_<95bGQJNOM5^Mebc\VZ6-H0NRB&g,2^9=Ae9
(&,(.4^E\K]:P-ZGJ;?+6D\-<5_2)&Ya&A?d6Y8_]9PfV5BIJ^Q2GV09O)M+b/R(
A\E^=)dO#6OFgC2QB=,N?(=Bf70Q7B](+N/82K@K=b,EN1,O9(00E+P@TadA3b.E
QdUW43PKQN0:IC2E0=\_XHOYDKfI]Y,R?6BaG&Y:fGc_0\R)947>[-Tf5>S,LNGd
@L^TR:e3IbcGN9SA,)_GR82QAVVE-A?/B2HNc/2a+aS]K,X\.S@5a;Rg;[M)+:.^
YLVEAW9H.HW](b,7R^];dc+JL>&?D@:c-A@]R4E[^8P:AR=T)R=[a0I0RO?3a\TZ
/<5<4J/WWBc=f].g[PSfVa[A5c<A@8/c^\;gLb>bTE(U\N.EY(6(^2=LD@a.OA>A
?DO=V;)/Fg]5DUP)V#FL-\U8Wf.0,,X#&G].RHNX\I>Qb#Q1:DX42I_XW/)^IUOF
TOK;,2UN-25Y<g9U:.a(TX^2@DbO.KBN?,LgY7WOI4INX5Sd=1-:3K?16;d9M9]X
84,LWeM92(#<EU]a62UOYJ76W):PFedI2Lc(WbNX?B<,e2(TYC2d/?b,+d_[^f&L
D,HVC5,L-]=O7<XOZ^&(F]]1.0a?81P;<<A5H\UEMI&>F-ET/.232-9A]?=gU/]]
:g:GXCFG\FNW[.;D.>gR_7LSaPcd_c4,3:6_R<LU<a;[CK>DPW1?RHR1Q^I0eDWJ
H==.(]A>^6c?1RG?8\Re3c?&<WL2)S/A/,LOVFe,[X7@(Z0E-(DD-159b<JJUCF2
L(B5F&EO,QZC9PV^1ROYNG-3PAfJe#3c),?(1PSDaH(7HSJ89WaI_c9a-K8Mf,(<
YK-&[W81[O<dG3;O)B1ULRK1ISF;/J\JQX3I_QFV@=@(]0/>\2+922NBOaM)AX3d
ER(,>;XW:LeXQN_DZ?.X7MI/4K5,/AAL8MaID,B?e4_3G4Y^cV8^PT1?UBAXE)#4
HTc?^E5:e4PP6dS]+dZOCB9N=94;BAM>Q[[>\WV9]1^OcC5VbXAODZ=.\7\]@;?7
0P;ZBObX;EJRGIQ6TJ<a0fba16LI@b657D2:U5cPP,B8[fD@UPD@+gb-9@)c)RKV
\\P^.c(D874\7S3d1M<XC/ZB_43ZM\-#cBC59&@KEd7K:HBDQ1W@GO76RH;EQEbF
9C.[Y/0Y37eBJ:\<;05SM\<QK[CWRP6M4,CZT;BE]D#H/A?f52d1NYRd^&cAEMCa
:QF3E:e(cf,EeS7PPa^W;EAOQLY00//aTb2e<^5-7HL(3L6M096<VOeX]^HcW5E1
g/J7.>?ZIBEUF6DYgO0@U/MKO)L/<=79WA/(-,GC4R31<RA0Y?0FcbB9CTN+_HY2
K]0TKbG+/Q;C7@9H4U1RV)fO[;==f6bCA6OPd;AeU>VIOd6VE<L/QT2A0H2CdBPC
2V0-IaO;I&E7R#+(Z/5;4M,YY0XaR,E[[O77(a)6gG4FG.X5C5#LdCgE,6TD&dQe
7M(gJXZQDSTR[]6_FQ=-Gd#bQ)@cD0VX^/LR;/eE1A.1P[(4&fZY-4PO7KgJ+@A^
@R8gHTc(@RdW]\K7TI44??&2QL_aR-Y;>J?-aOg(.Zae-I[>D2.b:_LZ96C#CdMW
G;:OZ@,]SK-]=Z/B:7CYIU00&J/_:;O,C,X,eEeLH3eXSMH/KQD0fYFO/+[DQKe5
[UEM-?>>]V^A_B:AKZ)b:)R@_P-<AGO8>X06T4-G/Z_0.(e4G5Z.#F>5_\^eaYD/
\?S?Fe-Wd+&-_^\KX1/gcVgV?HS[0.TD6?YBX]_Q).8JU8F6?:ZHMW,4Lc;@7342
?\#X5[Q,\4/U\C[C]X4.>O:<+MV.I=WW1(#c;R3]DP_N8[=dHC;Z)I]BQ=0;],DI
;W/(\+b71G,YW:.a@#[P;M#TC\M=7]HW?gOfGQ<?FZg.OCWb@-WSII>CaGV1M(X=
4^J\SNL#g,,Z]4@R,60b-?Z:/6Q[A^@>IW-:M^2X\]IIMT([O;,E)_f2A^/84JNI
(.4\@H]\Xcg2bH]5ZG&NFWA\JX>Y)aff,J@A&PMc2F]B<:f?29,TUXZb?A(d=\c4
eEN\CO0bO=>ONW11+EG^M3TC@(eE_+,LedK_A+.a)VGCF)JHaS?d(WUELBY+;M@9
3&<(HaBdfZC5UY@gXOe@5,:XP+I-\Ca^Z+T.SI=cg+e6P-_&]g7)aD)0EN94@Ac2
K&G3-dOMf-G?I&F&M_QG[]g\<??1UYP^\X<4MSX.)-B[I9JKO/1.AT^Q.VK=LAL3
TV]4+M0I?BQZHEJPYUE?9<_[YW;G[?W,[92ZOXJ#]>[>dFDTcIYPGgfU)325#/WX
R=^NWagJ-9)O<J\_G]4^eE,>AcHa7-8?-M<d+^C5[Hb\U>OOUc5V<M?aM&I[QdU=
@b&N-C8]K:ZT.61.WP7UW@.Ud(M^3:J+R:F3Q(eX+O)UJ4X+7GcKU6S3R,3^#M<R
O.[Z49PA\XY=ZBVK:&.7bC_[Z+g9[c_JO_OG&Q?K[>?_)(-\f<1=[YUb@B#PFQ5f
@HYga&:7:R3E@^\J[G8.0Q5,^-,AGNKS9/]X:;,;?(a:)AS.4S.9Y?LN-@([AJ8/
#=4<&f,IXg.@LcH][T^\1?SUY3bUc;]4:^:LI82_CK#c3_NN]>9c@?P2]Y-/VDW4
BcVd.<U\&#W^FH=UF?+@>)>UK.K:7NZAXW.XO^:BCC)W#NGV<RGC,986/9#LA9U;
MdEQeVF[-QLC>BN@EP/1L#ZPZ3egM[d5V\Ta[b=),@:F<YO3g(^OSB]de]JB4/b&
;:+gHL)bBT;HNA#1^=:D^.4TT[_7J>b@6Q[:O#c<@[Mgge_A-]F<.K637V<P:9Va
XX:2GBX4\O]LM8TE45DNMU9==7&#NbW_eZeg6WEA-I1CbZKX>2/?=<?29@^AN.8E
,.2fOFJ.8^Z+-61,Z;A_:(KaT.b)R1_g9/EQ6<.SZ_[Q]^=JAKeb]3BQBg2<A09G
N,&fe<6LHI#7abL&@>gNJR3Mgb[TLd&-YKHHZK4_6LSF]9L#=Y4C-ZSRb1?-.+[;
R?&,e8OL_+>^0YZ)0bV?QWcg-c=R36fBbU+6:0H/GdFWI<RfebXf4YS8g:S1;aT:
+BI>HDb:;;.cKN?D86XU1KZUZZUCc7MQ0>,-caX[;YC3T2WG8@-#Y3:<UKM>Z]S+
).W@6,VF;\160O>HF>D3XT7BU5>Ug-4]=H7H?KTYHY(8WHLDD(BAa]@K5E7d@H09
JXGR,KaP5fQ8JRUcMe[=+):&QL4].P)IN_67QP<^7ZM-@.ag:aU1b.&;6:c^\.JL
\UPC68N,Ac/7,PFH)G&^:6#]DWCb5YYd7\LX\6J4EW4HRMB/&@]0QZ-L>eV\=Wbd
R0?DH7_6JFD0Zg..O[]U3ZSKL7_<.:FQd90/_?ZTC>C&D,<(HIVB-E&.YMK&&/IJ
^/:dca^=V1fF)#TIX,SO=.;[<]4I4&SE;(YOKfZ9c:TBESQ;GDYY^U7:_?K1:4]Q
Ae@H(FOB9X=W^2@,a3dV@d/Oac7:[([dSHd<Fg3_gTQ-9g6?NF06(e7@T7P7_:95
_OYZ@f:C2I061J=F8WD+bc4@(-2LY1/;S=@P22f^VX(R;HZUdQLB>1236d?]PNAD
:H;bR#HAd::HYHYAZZD/^)C&GJ<+Tb_3672PeWE_a@GDeB-]&/I@9;#e=1:HLdW8
>(4SL#.1^79(68GaMd>9ASWYf>O:CdPE]A6;?be]Vf77?\)BI2E<Z<HFcNJ)5[>9
e3RE;?W[)M.NE5]Q7bJK9Y8J3>UM,Q@8?SI53DCM,:YZ7JDF6X@EOOG7Y;ZTI,]F
C81O0;HHcQIbcNZ5=D@QN-T]eC4_)U/GS5UXM7J7WeJ76fgg:.gff7_KLBgd45]Q
.R1HdH9@.6YSM)A=QO,>_a19dPW:D[Q08TW#;Yf)09JXF]D.EDEFZ1GX3^/:DgLG
]3N\WUPXd56YPgAFbMS;eF7(Lfd_de5@,/5/\SJC[(42JCb\>de;T@RZf>.gNLIA
a+0E4abVN\4Ba-4+JXV2>#&@fXIAB3[C[(.-W>[&\[O,e&GV]X@W:]cN/cN=2;4E
KI8[)OO.3J-@IV)Yb]L8]<M;ffL]9LGFK6I86e^);JC&[L@>QgcK>1.LN+H2E(Rc
TfgT\L]33bO<=gb^15c2SgcG(R#-d4X:/)WbI26&[/=_CL,@D>aP\-5C0RfO:4W+
4e9,23aP>G?2/P3c6(PQf1JG&-#WIe<&H4-M/,KX_/H-XNYVeA5D3\Tb=4T[,\c_
</H7](B,5NA\3R(JPL^>gPYV#TSA]g-1+;([EQ@9X+UG33][4Q8/&46#ZQQG@ff9
E\JQ@bZ.RY<:AMXQ.6NefB]>L;/c,c4T#3@(fd.<3<9+>BCUT5b-C-7b4>2UHJQS
=/RWBDQS?&--EUfB&fWCPg5?&g5LQf)(Q7,HB3IM,5\RXffWOSJVaNSC5_:KXVXF
JP5d#,)R&:bgTO/Xg]U/B5-DfS9bP/#+J9/.ZPZO_ZGGM;B-#0-DK^..c[TJc\^b
a^+HXV:@)HaC7F5UR,IPDAXX01M=c#IO-[N?XARI-;G/,^.L[U;Q5YbAf(\X;\39
/C4W.d(]TN&cZ9)<OZKeReV3C?=BHOOI&5@QT7c#,dYU=Y^XeF^J&K>:[,_KU)Ue
,N<\.e<&I8285TWg3Q1HDcO,d8dRNX=O.VT6C]8TaL6<dSNHYWSL;1+COTLTZ94K
D^>S--O=5MObLg0[4cPfN9L3d/O\88V:SOc]FC&UKGL<?T/L\TB2](+X^Pg3eGOe
(I2VcaQ)g+?EbQ6#U\dZ0SagUQ?IMS/F>RTHUZf=Z&>2TVKf\K]dZ)5>,,JWD0Da
aOESIV?=6fgBd8/bB8.fM(Q1L8(I@KGX8QS:65e0QU[+YaF&[fT3N04b:b(5g1_>
4ML^<Q)HY:A5+TZ+\9c3#e3[IQ=N>d2T-&PN+geaTYM]#,b0PL]R<6^2L8;1DD0/
S[IUUXM;4J)Y#Dg]13):gHHE;BK9S2gTe^K-bW()#ZVG&C986R>+0HPKRO,].UZB
3LL#1<(N4\e4OOB__HXM9QY2]cW\&[[]S,g+E7VLR-([>fTFAZ96Dd.GUBLRV15b
JX=KZcbPZdbY)1.IB0a[06GdLQ<Ka5Of7EcG5W>,7c[@)d:9G[JQd32)H3NBQ-K_
aZ7IYU=NX?CbZSD-]XP=77HFCA]<WT=W,?2Q8a>X-dKc5Q#S<PWY4GJY\PY>LKcH
gFd6P-La@2VQ;E#&1Y#cU?7]C7+IQ<e-EWZVYb0_B?75\FUJdX8B2>FQ&NS@Z2U2
/1-];8gf&F]L]\Z63\IZ,PXIZW9V64XKOSO&N.LKG@c09?6IWHffSLJ4=H6<JW)f
.c;)N.T0H8J,12:dD3TY7U8[dY(aYA^LP+PK5EEfNYG,PS=0VI0?2J[bNG4/5@PT
FN.U>/1/QUW0HA04UX_@M/[+DU-^<5QSBVZ5>_]_RK\SV7b?D->eb#.ZDW2-XfG1
Bd9X4:gA1bHAXO5^,U8GI6G0TT7DP70?eHY2G\O)gaJN#4TCL.?,B6d\T?\+04/V
FYX,JFICDKALUO=;QY<:7HU&78)(-C]N;G;CB:R@\cHVX06UX2bWa\-:D]4M2<FE
H1a47;2Z4S-)cK;N^M2E#MAb^c+G+d:@5CDBR.3R)=84TQ\4((<_@f1JC((Obc4H
G.EYY3gO+>M-L&c^E]FLDg,G6CD:-.YFAeNc9@JI2d4T:99b.>Sb#9PGC2QaUg/e
Je<>+CE8\11U(:0I&&\JVWFG5W(W(U@-#83JeUFL<@^>Ae@QI\(Z+:C]7E\ZJRSX
,+D^dQMWB,dFW@Gc77,\N=f[]=0E5MgF:71[&;VO[>,B[D?=W-@A+aG@^1-M(8A@
?&2>NCOP,BAc2V5Q[9]042?f9cXB3\A8P0?KEY(R(QY61R7=TV@-(aSY.,N?,]\N
4?E[S03:C0g8#HG\.ELV?[>]]5fAH^(=8fE#2;))?W2Z2ZYIVV@>:ILGb@P_YM1T
Ff3e9D3<:OUdHPQK0L^#c::@MeM(W0N24&YWX6W5f;19-+[+92+1>@S/QdD52Z>=
JY_U+\MID@OUAX5T72EB>R0+Ia5KA&G5YU([3[X?a.dF,LHL2>OH/W8dXBFNg7PP
.I8A@8RbHCOU<2J/T3RA1D:VW&S@W])f]BXX_E6c2KRT#_9RZ#U4H&b)C^BI)YAL
@g1D4<.a-ZL>Ag\BbZe4]>b#2FA_F-YBHK&S=AeV;J0(f]:G.9fG_I=W9D7;RV,4
JgGEFH/?BCa>W(]T+WB[-Rg&:/=[5\M[;JIEcN8,#Y>fBR.NH0ZYF@c63?D#LP<U
3bf9/Gg&#bg67D.eA]U-68[G&KYO<cUT12J3@NPQD0BCLT.D>P1Z[[C#3R]Q=TPa
Y.4BZCde---<SgQ9^RgM2?(Ne:a-e>dW-aADf&\b[]EF5N^dAC3N6IAfCbMg]:&>
OI3J[H^^:UK=Rd7N2Z;[_)Q;D>\9@:bG1b^PCG4.=DISG/2b<Cf]@;[LKR(RU/?4
c(,_6XE3W-Xf=,,/5,[I>07X_PY?(B[-@)8V#,O:A(Aa_aG4)2Y7WQ<]aK;89:J.
_-)FC0[28?,?W5D-baWGWg3;ZD<-=_LZJ839gZB0[X4=EfREbPY1+QV0a)2?>XSE
?Ka8IDOX__;)E4D<YT&2FgBcIFUFQB[YG(BJ_]@H&8-F_f1e^G0Y<+E>=@gW=;b1
-B0.E0\7C_[&^@)(&/6&@7KQH5]1)C_Xeae6<9Y[AX2ZVXOFH83U2YKPFB<#ae#G
U2G:R]RMeN/VeJc]MBW;ff9M2\3/7?,S2Pa8(N0121=KOI)KGO7=E9W\&26a>3DK
EN)?Z91a/f+2aV:=)>ZIAQ/HV8D[4,8Kg?fUTS2G(d06R\22]ZX6W_8)).MM2(@(
^&WgX^/@G;EU@a<+--JEN7b:)-+(^);f5>D^.I1CZB)MXD19c0I#JRKQ&=+@RY#P
1>@71eTJ29I4eMO?(bOZC9J9.)CE_GO<V+0?WU4d4G1^A?B8&/=fPT(X3W/f;H8^
:D/LU=EfJC<e\dHK#9PecW?WKVD)S0S:b33Y?/JUSUK@T4.MN&[WOZ_,CJ6SS[Ig
2B7^M2TCdDD&JNb##2]Z>Z:2fMI-BH:2#P9eeJd40B7NF-J:6e:KQ&fL;dG^2FC&
A0QZ^RDSOY^c04Q^a/PXG+W+5+YEV535g:O)@5.HfO[F\:Z<dgbTgUAbB0.dMF0D
I83KK5\6]^)IK]QNY4geTX>\09BQH.[.@NXBf>7QD?f>7O;-WHSC>X.LK&^?0>8S
1M8Ed.(L8PYTWN.dM56:@N#(QM84_X=+VPHD2<Q?Y\H>CdDDZ6LC1XX9?Z8EbFdR
?aD<[2Wa3&S:D^(-56>W8V\S.LTROe2g.Mf0?6)I.U@#cY-2cT1e;#2[#KA\bY0R
abK2f^g;J1ZNRR;#\;ZM91be2eN#f28T1D&SEPI,W_QR&a-f+1R(J@M[IFC68>E<
?#J_C>JgE9d0CJe;3.;5N[RG.cMXW\-P+cGdH?EBD>^Y#Q#afLC#&:LIaM#J7@[4
Ig?>#dBUUY8]ce;P>/IB_fA<+8;:9TK\+aP4>,OW.AONfK2,?>fJ1WA\CI6I8WK)
A4],RY\N84agNFDV&8dJ6&gc#,;=dP#Z;[H:2Ke3c;Ec^^UeVJVY;.M_W^X6f-X?
O&IgEgS77HX6I>N7H],_:(a.RKKT1Q4LQ647GDF64[@1+#N,:;.)EfBgR4;Z/,-2
W#OOQ6@G;968]dfBL6._KUUQ?M4bTXDdX>1(/8./TPX_T=89DgA&.1WXP9JVV^c;
L.<VRK[-;HES06D)-STP^Y,_VC(4\]+<S7=Ce,fLfC4@2-XYR(_&3?,).>N=D2F?
VFR[7&[^10A:#Ld20BAIB3Ca&GKZ71.^_P-YdY2\EZOE-CVS2D4L3F#V/+W(RK>[
.aP<@ggPRJa.E;:R2-J7@?:AE3VU[32.4GBa0Q])UQbPRQC1-7fS(9ONPKVFfPXN
/C>U^?;g?OI<L\UT+=]YLa><KYXccYOaQ674f\C=^9T6Qg3Q=a\3M8.&NE&3309@
\&NKE@Q);8/83OGF_e/;&-)R4S-LGB;b<&W<8K?4TZNOPe_?^f0C(YSb,5)O##>0
LHK-<Q8K^be-WOTZ8WRCZ+-?&aO9DRQ]>-RG,J4:B6PM0^<b.Q\,H+bW)9Xe61BR
H8M5>XSLD]<7ZX]A]KYWD)b29cYX>NE/H&G;S@D@XI.e\/]HG2WT_+e]/\&=]HEO
(XdaR^2XVV1H=>4BFNQ9f#ab1RLRKW?1H?bSa&E&\\ESc-(3Wg8/V2deZQT\g,+a
E3gLS?ATZOTV/QIggW))[[/)D2?G,?b(R>\7YBS@;_<g_PJDZe\-dKUA,Lgf8,JF
?QCW[[eGRD=f6SWS:1c+fI>YURH5A:H9NZ+<Z2@7XINO9_c1)eIgZ<.,2RQK:;bG
\0L5ebB:?2JE36(1BF,BOg148cSHJ?Lf[#G[Z1SHFTTXMK/,4)0+S?<;T]B=_LZ-
XcQ6?&eea>IeId]OGH^]JESV)>6]4;(/872LfY(V6;Q8VH74]H-]EJ0K]c6I[dc]
>[b_/D@08:CNeK5N[25?_c@>LY:d6OLPS1HFO6IKH)FESAE2SX3N78SEK3#R79<J
\6Z@J,eFJE^?L(D=EbH74T(d=(3XST13//+-dB/K+G8H)/I2(HA_46G+4B^38?#d
(T&DE180=PT+D(GL(M>KSY^;/8BaS<K12T892e2X4c6V<aU=C=_U#bg7LU]_SUWf
I).P]&752][S_.Z3QT:E6DFT:gW5)B:RI\70PGH=^Ne;;JVA\@]I-G[K-M=9L7H1
_#MB:^EP20K#+Q#=H?O0VY@Y4I9X375S@X5XE_&GODZC&V)(X^RPbgJdQCe>eZF1
9J\<.N_ecacDQ-64#WZSL:L<;1UcTFPXbR+.^>NL:I6-,WF>PD:+,:+>8.)<]1#f
9ZKf56VCKbJc=^F(a33aO2<F\bEgKfXLdUf7+\IHMbF:T1&&f#JN/CRZGcYe(K/Y
6gBUPaD9ZDI=-N&Y+35VMd->1Y^SL3+b3)2B>(@V#H75T9]GPB\[fA65eAA&eK8.
G,:]\O\/@W0?K)bLZU#,J9OecH4/f>gMU2ZXbO@:TQGM&<fQ#N40H?6?GY\gK\BD
SA94GeI,b#cb1WV^7RY9DV?(SM,QNfdBY9O+8M36XAVHL^Y=PV<R_7>K2<B>1O0(
@#211CK2EE:g=\I0<9S6g:S[^YZg@<-Xf,f1R-BN,gQZ2-SU,FV<FV/:BfE(UUK.
KfMb=->69N@F>b,7I&=<:KN;,NT[dU@O+?QL9LaVW_AD5b=,UK^&a2(19(CaR^UN
0W2<a:HR(9\AU5>\OMTLTXD]2Ab,CVA=Y[.I(C94\CNUeMf0-CaU?=QH&Id4FX[.
;&4C@Y+MDN5/Q@7CG/Q,f8d&eYf\2A:MY\VD:Q#8AO+3]YeK-@PFW98.[O)K4U5C
ag<1WXVB[dMN,dTF7^PD#_3IU5>a^==81&TVHP](N=.SB.#O)X@FR9EOc9g)>^df
ZH7#^D0Sg9=V^@T2;]_ZEdCGA7I_f(V4[4>1Id9P<A+S@f5.KcP6\SE1O:2/05YG
C,=1b>+G7dIR+[3D4f?.VZ[)ea:9]Yc68f=YOVYQ]&R9g299AR]MRD25KN.10?T+
6Mg]5IP[U<=D:8fX^5cRC9gT,.W+R6J^N00?/:6EC^7^-TFWfP=5M:DJ\P36W/eZ
d(_a32\HE);a1Q2=O4MVS)gB^gcB_I;4cVIWBS10=/gE@F)^FdI_7D#S]I14^FB&
M#<26>b)6GcD(RgNFH7<4\+X()R16eHN;>aNBK>A-(.4)P[SZ>CN;P8O?<FdRd#]
]GK.0PONB_LE10YEB+3MZ))I;TNa04A;UH4[3PA1QLgOX&[HXA(aV:f]48@7Id_V
MSgVC?6ePH<(NWK4URI>:LFE108bgb<[^>5#[_X0)&^EY/FZR^+VW,]PQK[X3IA/
T#eR3F5I^+T[YQNVXKMVJ7KM:^f>;3#cAGfMQ1-AG?+;aYW\FI+ET\PA@+F<?<8N
?&[017fG9ZbNMd>&,Q;RF:T_:J?_DJf:DKXeA[=bT4?FId:RF4</H=#.+>I4A\14
7.#]@(?2;#WB=(f..d^VM<W5Y/d8bS(7T9dQdaF1P[.P:>(f&TZFgXW;Wf^-Q:FF
85?-[eDC.fa+CNIA3JDT:TU8dF7LdLa0I\^V.,-;?7K@(7TfY@-G_L&M\9907)EC
gcQ8]=AA0K)SEP7c,TRFG+EW5(1d,?Ma&M&d-/f#228ZDVfA3d2U6b=9=aMWW#<+
#VF.FIDB=<&RN-Z7ab8f^^\ZD^0)UVU<L,/(KUR9>/O55feEHD_#6)Ib\HPg,2GF
TB14[3>VfYQQ0:V^fTA1GM21L[O&)9UI0N5d:EBS:X?YCEc-EMNg82H\GXF^[(3Z
=1FB=U#OSRXR502/IM(_g&c?-[&8c\JF<K9;TCd:S2QZ&4(#P=d]6-,bCN#D?&ZH
6:JYCc&LZRR;\BI]ZSXa/OJ)=@QcRDU6LLAN/0+3)bfB@<CHTEb5L@V0-5LE5Z9(
1H6?U7fe0OFD)Nb.ec3)57SR:)89#7RA@PUd[E.HW[]G&#AGdM8E?65QP0)[^^I;
\].),F[c2?VKY1C9C<F.71:@]dQ]VH>XI/T#ST5D@_#8VCZLLT4f7-5BWI3XDS5e
1ZTCCLTA?39N7RZ1c7-&URA4@A/dMQ@;f\WICIg>3;?FDJB3J+B?8g+:T[41TLPL
JLWaRdZ40a8],V)718@23?KW.IRNB4?^1<a0YF.T_&R8JdWf#(c73AG&W=NOY3?/
eX6S5g:;9fM77OXCJ55O;e1cac09fNB5g;J14T.4XHAE7F5NC3Zb@(LXZcdfYR>)
dL#,N5D:FE<W&:bBa:HMKG>P7H&@[=7D2_Af[+;>;1IJa?QfD>R.VDIKZ(RHSXSb
#V5(Ie3[V36Xa#TaZDHY^AYJAcWV^F]@d&8Sb+O)2[2OA=?8QbPc]78??Y>P1Oe(
P[?g1I:Z(867I37f_=<E=I0,DbbNC<FG0dWU[f<HWEWY_2305@PRY[b2EXDJgDE#
.E>1:;U?.IYS)0VVU?CBXEgd6RJBM]-M)FMgGQY\Q;/S,S1,W8C?=BW2AM]c^ZV5
,=X<?gV_9F#f7X_3?.C@fGH\?cZ<8THKY6G1+>L]R@g_9?G0V=Rfc41K:a/.9EK?
.BZdJ&f<TT;;8JDG:T<M1SFJ2XV(@^:NOJ^X,Q&,K46_ef[8Lg9[1@_AaM).35_<
ML<<I:?M/JI/_:0HN>86d(]6=6/2^eRFN8bR1[ER^IbZJ6C_,(2V]ZT_=76BALB]
FW=,VR=ZDCZC1Le(YAT58E5Q)LKNMgH(U;aN,=eA6NFI-aML#(-P+41W;^gHX/_(
HBZ^S0AJ=M][.#3cZO5G&Ce(>MVO0<TSOJ+17-J^+/ZWRN69,gdG&3_[IKRWS,WE
Ha=@#dZ@AO]W>2U]4H2LV5CI85e[FLOf7^,>e5bV]FTI@K6Ie=1=g0I4,WYba,HH
-A(<H7,W2ZQeUfZC3MCS\U?c.=?@WfD<5I/DEZ58>J=WEJgG0^7U^HNaa60=Ca)2
DQe,a;@D4,AY4MB@52.)&+b:eVM/IHD&+@13X(;G;d=KG8WYOB>5F[-(O4B/Q_,?
:4X4_G,=8976:=W4bV[DVMI=>FG\#@A@SNRQ3>c&&W5P&c_JDX:C24TG0[;=bGOV
5@#Y.cJC@BCG+J(1N9dEH4fY6ON#19HTK4KSN/NE6aLJ1+@_I,IAG]?Q1Gg(g9d)
P47NC)7(UF4de7eDZ?g_,R#?D\<E3Q[IPLZLgd0&_EL4YQ\K_;=6T,ecSSdb#&I.
eEf(?NT1D2Z/=N1ZGITgaT.ZTY_NU4KTFP8I8aX&=X@+M[93#4MFO?=)[8C9>ZHa
OT\-:2+99SP>E2FY<c9^W>6@O2057+M:XdZ71gS.?CQdYICH753V>))(.645B+C^
->G?8HKDBUCgC0DDG2c+FH>WM?W\eXM&HWV\M=8?UcNSK]9P<<GJAVY[/R1L/CZI
PQc/12X,KH7NU#Pa7JBRVBY?caP.YPfFEF/]F&fcBMTCGO<d/;g=S@agI#U(UdFU
P4[c@\93<3/9+@NR.DWfV5]CE7(9G)()&O9cCJ,7EeF=gW9:Y#<HAE[==TcJa8QG
DH]b9#a6.gb[Fa_D6ELXc1Q_X./ZdA[ZA;?(XB33/R3;<JBY2c:N8M^M^MW3#<.:
.,+eJ&?27AZ4\2.0LS=bWG1.gf?\\:=738-NM7GV@5=.WC8T1UF6:3^)&eZUKF/Q
(LGdO7(XE+Wa=.)9H?60V1QUR9LK?4Ff<JN>&7aUR_B=V=>;>Y@?dHYF\F4[;U2[
S=.7QL,Y@KSO,c6G(e2:WB#P1)0H:Zbea_QA/cK)f=Kcc(Ac=3<eHX^5c)1T2]K]
NL=]>9<dMKK,N@/0B9D1bNLE^#KgYZa-P^\U_V<ZM9-a=FS/;02/&GD/9S3X-ZI<
cI+d6#Zf<[bWI7U;MMSKKP07E]g/]@N&)dSJ,DSIW#XIP=DLdN-J&#CB^./5aL(S
14PWPg.J(LbabN&@-gMO#4S3b5<1B>/4.#C6e=IHKeU#+MNbUGRJ=1ZZ9/A;S@><
>70>:Y(6N7R-7W5G)>P:2/T@XK]+9aPI3>P>(BW5R7gY-OD)0&[AS<TC/ZA77K>O
a(0/M2>0f1/f>;:)-c;_BCAB-]XDb/))8G(2:HT?g4CcfNP,.;C6+T48)QPe-S)d
Ta(?8ZMcSP/-0M6_3#P(@83:&d@36bF;ad3&U(W_5afbCg7XWO6ENJ=_MT?A85HT
\4edHK]?]JR32^/?12LGRHM2/TV.82/f#4./_@d)9NfB=?1&?HBAO8-1AF1RA0M?
U5IfD9JY9aVSN)c5aJ[d:E1RA,5Y]?a6O74d]JJS0a.5>WRBH<&a?:?[?JA:]g4_
2,MAdIYFg:HBC\<;BaH:<cVC>HF;,Ad/&N4JQ1?;C/Ue<dGd=2B.F<a=+fFBLXX(
W5DJ0)1N/DY;Tb3XJLaZ1=[BWTPM=KUIS1?/Y/b+&G65,]^Bc9Qf2=UOcH:C7G(U
QR.,cLcN(,e]1XH]/Q6bSPg+AXQg4\:6;)Pcf:S?.::93]#cWP,2#Z1>N1ffM/2_
.#HN/JS-c)DWN6)HHe3Y1=WTUX&F^-O-VLO4b:0@O6;GJ1A^XE_ea@]aGG@QgAJ;
[A[DP+<:YNAJ\CQ[9)Bb36D:&;e_^QRM)^[;+-TTgc5b/P5bOA,[OL3@cVDT8TVb
5DXQfP#L(>AC#I>>]5aG9>SD23TP&H8O9OR\]^OO2f<YbW_#(<;JR4.@>@]8d&_8
PFg86=HeecfXc1\:XA&FF4;]R[9a5?0.P36:FbF8#:,,VO5QT./\L_KCGT(P]])X
QRI+4#0]W5<>5JZS^0+]874VYcgKABce2MF)1VD<Y,1KbeJVUQ<&V>-(V:;;Ag+L
NJ)R&79)09.BR-U^Ee#G:OR(C^_cH8b[Z\SC&8[34R6Y=,a<T;(7M@YIH9/P&G;+
[W:X1K>eQ=3Ec]^KRX_GN=OaD^4\N\d);gRJ_F-#5&[#\)MRF7[[N_V(7=T>gI]6
9S1fP5[_MG7DQL)e?OT?ZVSE>cWD]SbJVD<?bfb8^JB.9,g<=NW8XIb<LZ>;3<\1
ca8#3PR3PG-3#gTG]d:bc?E(fU22G1Ie_152=<\)6LRDZA&3YQ=5=5I3)cHD\Q>E
(Hc[1ZG45;N<I-V-4QO55?W8\gE6TK+U+AOT_bGO:EHXcB;IY:0:XJI6.+?\YK34
5?10fG(\S+&>@5+.?00]2FKe>9=;\,8;(IO;</P9KB=R>g]g)bD:+cA513D[0EK=
VKUB\LQcH0d)\\J@?U)<BJfLG^JQ0?@<W.1BE5C6VO@G]L?dg_R=<U^d3S>J\KbR
<1T?>eDABUN;-7;O8V=fS7YHZ.OaV00VPFN3;5C8eM&54/AHa3C?L=E6-a6ObL9<
acZX[_aF?/-\L@B(;#2@0Q0c:W\g>+,dVQ&OcTeb44;N&7(XdH,/7B5#6>EBS8=8
G)-2PGU:#7D@L-aW,Z@RF?-M@F05O7[;O0+c-YGA9LS&]E+:.IM_70Jbe2E48A9.
755R@?ZML4.WGKM_KO7GC;@X6=c7fJ.?g^W[M&^8K)77>B6/fP/N/^RRK)?1&#0U
Q9GQ?-5#-bbSDdHB>Vf_LW>a;ODDC.[;CCRU/&FG44<P&E8[+dNRKd,eag(OFSN-
6#=#4^WCV0Q),D(NQ4Z@8@0IVL:f<3G[5.3<G/X.H2/7S\;>W59QZ4,<16\L#M+_
CT@[BEP.0ZMS+JdJI]eY].G/SHB7c^T<K=WC,\V-JX3)Pd\ASC8^VgY>YY-T?[a&
OI.V1^FFLBOW#-fWSKQK/-XFVE<6FYWaDf:1HGF\;RDLMA:P-0F#-][IX3MR6)<+
(#<28XQUP8WG_7:I;:6CHQ3;g)CZ4OU\=?PgT,c^B?_=[@HO;X?-5<E+9?WeGUG,
4g]A7X0DMX-W13U1_XUAY^@]&UE]Q/#,K.fSf-:CEZ)F?4d8\(W28fE5eN<GXQ-9
<R;EHa80:g857dSE:S+5KL>Y#@S3=,Re9U&ZQ=QbKZSdeedFcXLBXeXEY-VWc.W&
cVP+#&7;F.PDfH3A<#e]PP1gHaL)6W=Wd11#=&0:LI3[]/>TEK\G8TKQ):d9f(KA
:S?ABeC_@,8Je(SF6@/QC#NWA(<[IJ3a0SN3()5,W],0=7a_L:gZgbZ+U3_>Y]BN
AUP8Y?2^QJ)fGfRUdY\JRYBX<fN94_ZSUEY7,Ub9BM=J@_27C\+?U.g;K(EE6T-7
@;S78]CE(\^_731UR9U\=[[;GX^<3cecL?5EcQG5U<DI,6bWY[O,>/.eV/;R/OIG
VebgZ1Nc0X3Zc#>=QKDHFeU&cHF4<K)2#+3)^M#F7_VHE0>J<_]IYPK((II[W/7b
@^KU<W8VGP7J_,8a;dDC_84_9FRB_Zd-/+_XOU_b16RG]f9_2ZI2JINQfb\eLY&\
4#<Q07f6>/aS.F^\_L&Ab>a()/#?419-/Mdc&T_Z6c0@;DF/5GaZ3=51cb1;aU==
F?3(?-;TY@67+PP?C/E_>?)LUZ5O:+e93b;LB_+T=C(8M1IHOeJe3S[>Q?#^8?R;
1VN9Z[@8aPI@N6^]B)ZEf>SWC@-BgC7X5@U;?a>U[;]EN@52a+VYB,b51P6HY(]@
O._RPb4Q+]5HCY8H7#>U)K47EVBQ6GbeOXfO;+bfI/Z&,<0B@VdZ47]Y-LKEDN1e
3=3W?(]HQ4>bW3/+dS2R>V-R6/&>FWdUMbO9I<0.McKaW:JX_?)&[<[]ZITe;>f-
.Cf&BCF383NS6O+gFXZ&f(8Pd-gW=?I)HN8X6GE-^?#3VKO&C=LWW9L^BMCFK83[
3Y[CZROcLd:<dH9:)Qc7Y1Jg\LaNe]P@H4<Ma>VS2+R,J[H5G1Sc/WJ-76/==@YU
SbgJ3/TB3@WANQVC&EZASJ]U3N3(Y7Ta<2]#^@;e+_c&L+VVdRWD=XZZ<6T^gCJ,
E0aME/VJY9#DAD8Of5&1Q3RLZ[M6(_cL:e;_G.#\O,9^>7PCGc?fK>?WE2[d3HJ5
+LR&D,/L7:GU\R9P=#gea)APA_MI52@KHHR0^ERDDUL9V3;eg:ZL@1dV[CFa>E+\
E;(AWMOfYQ8C9&+/1FM]1BE1?cWXQD3TKES5X.5C]XYUf9S&XY8D>VW@L>_A9[5D
49#A=J>;DYMQ/RaQ\/[c>e1a[:+>/eQ^+G[\AI+Tb;Df+XACV?RWHZ=3UHW>9_=-
ZC+80bg6#&Q4-3gMVZQ5)WcKdcQ\N[021G-0TL)WgaLH,1C<fOINJ/G?5SSI>G.[
[)dUe^IVaJ=+Y=F5B9F?<N>,R)3<9=OfP8SY>N,01E_2H<+_-85R0YV+9+][e_RZ
7a^eBK(RRW<0,5WI^>@N+@<6>H8EL/#+]LD\YU+B&^VD-PaS)RY.LbQfHJ7/?A<[
#IJ4YM7\_D-9H\\Z3EY>3E:SRJAE^e]8VN]c=BQ)]bVeV5ZRd[^H[=&2?Wc7I5I1
X.UcJZ<#eYNXI/D@.bAEH(R]O\B.4QN(ZWD&F#b0X=82OJJeXL?5@Eeaa49T@@19
NYU_PUdPRbV&A38:J8M8T[O4Y4c64&</:[@Re?0Z=4F9^;7HdA(WNgJ^,.MCKG^3
XOML,/=A7c:QLRP;/^L9R=Q^-c;S^IQ4gJ8B)(F+]0?TER\TW4bDaUaBC6\\#?.&
DFf8@[\HPRXILUJ0RDU0Z1B5@^b+((P_\/5R162WZFMIeIVK.DCBKQU^H<dLeSGc
Y]cLfH,&LI;,5+SVAJf/+#:G^6eMS@AYMX=e+G1gL#6<[B#]495b,D8g>)-(\U&e
=E#(d4(GU_PX=(__NfG)bJ9BgAY<B3;g;X]16\7#8e;fU#(\#PM4)HUGHeTe#b[2
U4XQd580/S6X_9LP&aCbg59Q?U)/gQ_ZL5:&MOPAWKTDBFINL[cUU1S49AceWM=A
3I:AT?,D\beH4E@+PaD=/R_^NA_4:;SOVDM1_gJ0=&>C_2CO#T7cfW?Oed,gIS6K
:@BQ)^eEJ6/;F)L8e6F=DEUPAC)791/&(eIYM4F2KGJ.M+#_EL:[H27B_fSSYLdB
=-M]RP:bX9XB#TXeaB/QIgN4)?d(R)fc#LV,gbZEEdD&PgSIE[F0fX-R34HVUFS^
4V7T4\<Ma;95(Y.+W-#a2E0M.4J<#SQ]0D7+.2KDW@LJ;22WgYU^-]6__dTFDY8,
Eb:V:>[T)f<O^LR87HSW4XK)fV1L6?3UKI-+I7][b,4SdZ(KN=3K/]K[1<(=Y/Y,
2RBZJS;2-_VM.O]O5;/\^+L9g=f0029(RFdA6HfY;OISQW4)W,KaV>+=G+I5Ff^6
_YI<Cb1S1>JQ;1:.bG-@eW9g)/?619FM=)X7F&&Z?0K(C1EXARH[LFSBAK#D^7e+
^bHaK0#G^@.@b=HPS>UMgDT424<7Z38dXM;L73;OC@G^NR4G+>U@][d.W]g7UScc
MT-WMccNT)NU>:FAPTCO/#baKIT0E:_1B,XV.M#LC7-eg,CAGf=5998<MSMLbYSF
YW3,;EOHP@#+_@HH;<XM[V<VNc92W_\#B-N+5A=[QS8HEO[3)6JIQbdJ_G9.3S?0
V<fOW^QE_COG57X-#LSH-aXS.C2Q9cR<R55gWAIN=8C\FO9_S;-&)JA9.&+b^SSO
OXPL,U6>+XJSQce3La./Vb>?)JVR2)F82QG-=3QM6L^A#GD@\4c^<\HS&P-QN7B_
J0-H\FER(:QdA[:dR3=X=Y?ROX,K/&I)3^/=PV4)C@JFg9CIBE4B]W>c+(_-B,_A
,/Fc6-^=c-_@DeGBB.VWKX6PN>^c?BM(4Cc2G(#C_B,?b?^^GBQ+ADTTIad6N0Yf
SJMb,,4W,-c-AF\#5YI8Fa@5:-YK@8fJ=:@.DQa.74#ULOJfW>5V_V)X6aaXWEN4
SfM7BC7N]eS-c#8[;NR/\8GAMCZQWW[S+]ZJ?f938Ea5+2/Z#3;-5PQ)MVL&40[W
g@AT&6/dW^WI]23I#f&K2\CC6Od0#AT)egb/808<HE=CcVb3CKT6.SNXV5/Q)Ba(
]+(@g#U0IN[1IN;MV//++8U6f<34N<S#-B^fV<I[JTe5Vg=W7HKPPTc-Dd5Gb\EN
\MYO:K-9dVRDISI_3E)H8K)@7?Qg0)P38\E39D3&aGCU_g1DP5TAJ[b\DOa49>WI
ICJW167D4TKa&[2bZEFYd#U^DabE.R)WT@A2:FO066]bIC][IN^:WcG2LQRACSLD
N9IUH.6^MJ0NWbCc)M2PgMH(@aF1#,9&E_B-\Rc+(L5C]M[,I\E_Sc-:Q4S<21L?
9IPXI#-BbD,_[UO4VUG0R.HA4;Yf5SM:+g.8cdZ094I,cC[HfcE^,,_1Z]3^<60P
aL3GG@[D)I<F_Le9a7SA]He?D+UR1]aIFFVD&G^&G7-;=)]]D2M0>A7P^DdK5IEc
Q66/S[ZD<H\M1aUdDDJJAP/WA@/&FR9UR=DNBL2:)Ac-(Y;&e9FKSJNY@HQ@/^SL
SHF8<ZGTCQYG+B3P\[a7LP1-]?(0N^):])+K4g2CPZU[+G?8(S:/[45)EE7B)UR=
;.[>Bf]L+::b/Q:Z808OO\&3(3.-,0cNC-;WBAYL^NKcL6B;ePV[fLE+&V?HT8B1
b/b/^I^?IRXN/S]V0C-M5e-8SE65]JgNRb=?3?ZJYELEJ+cD__aNN0NN.@9BE(<L
X,5?HR6I7cORE\6XD:<Q>@[@[S[BDga2)KH>N=MZ^HeB_-)W]P)UX.VISG3_K:K1
d_)D[60aKaHa5X3g4D(P[8\c_RMbXC?fM#RN_,S9,\7d4T#+\,1Ga/-KTB5B?.a@
fP=02V#\I&>bE9=]L@A)cNX)WYPaC9M?X5cDP^BIQafM:XGX;+4TD1dB@H+.INLB
^?&\5N=,d22T>?UX^gUPUcT=e(/^0[)0-cP,R(6Z5J,f-K84#790(Q74ZWX+6894
0&R&W94S(DLHCM_>-+<1MV+5c>:UKDbM&Y06IVR>e9380fe5c8I7^C-VR>cWE+;3
PFQFGCEUDBMZePBd(?FO2fcc:W979]+>CN^K@5Lf:U#@dI@LQA^9g6M??Y?A&<M;
.+Q(K(&(V]A^SC.<c4.8V,HZDY5E2Hb7>BRN)WZ;\3,A]S_W8-Z:,7/.Q\S4UD__
dSWG5V5=cL22C+/K?:F2;.ad:Z+#d[DXFZRaE\:c3B=,STPG<EL1X-Y]&:XJQ^Q2
9:CS,7Pg<W<9MKXJ(>QD#GRB86PYS6eD[OM/6H59XN,XS(Y#(O+JWN1N^2W\&BU6
[-c.Ca4f3+Vc(&,M<cH@\VK#R.:9HE/>];G#JP+Q,<1D>B0W^.0cG([.T9^1Y\D:
^BWeL(BHP,?W49EV9<:A86R/-,Q<edKgQQIH)]M&AE,RA6+A3:a)_+SUVJ@c=?Ua
c-VXf<0O(FU9cTBV],+@OcW]Tf.2PeMX]@\=;gGZIEAG<9GEOGS&g4N7<(8BK03[
OVS(_72U=AMACSEd=1M[b\+@-,>SQ3V2MO.POa,3;>C:DYVW_Qg4>A/<+>BI5?T^
XePDg;g^_92]ace)H)9JB[bOd@C[X7AAVR8\@^)EYV0(AESDM:a9E=^]P/HWY_P)
-<Y>-FWTA89<F9EV]L]G0/8&FdK8/2bcOR@HgQN<P;9R+,_@Y]9dUVFe8WcE)<35
a(9_9DW(8,V,V)@@Z=Z.cY[_[;=^aa8#[S&9A9.AVH2?V+AA96(AOVIPRE31.]V>
0W/4,U,gTD,[gXbc8gCGTZa.\,5Z3Afb.+J7SC4ba#G9L0==aR:=[TO0Ib5DQES<
aW6RgY4[L0E,38)ZB/SKN-NG.K:VDV_)#L\D##[6T8aLNcBH2<BB)SNVeE\)Q982
NM,S01cW,MdGcM^U9;1TCW_U=3K9bFAHP-1@5FV;GE6>gK?VH(&@I&HK^Ke=#NeB
7B;C463gaR;8d],g?\OO_Z[1-B(B(5[g=7F8FQIQ:T^D@Q2QEC24F.8<Af3-<CeE
ea\3?BQ_<W6Aa<.JCf+-,e;PPE66_,5L>gc.&;,PWY]7BBEBFD=)B)&:OYaKWBa\
;L(aL+=@YSP-Kg0H1>[TG.GM^8.GD?#:D)@[c]d8NXKOU[0BAc(DZ=cQ:W+;NJaV
Kef6f#-M?GT7-CA6g-P=PIF+1P7d8H[c,OR^/B?(E?51DZRBK<ZUU/+OX_\CRR0_
J#Gb,^GKT+G:R&-d3^9=aU=/XV34T5(LV4JK(_O57H:RM1QS4XbE@[PEZE3_b)Y0
SI34+9=aIgOAX<fe\Zg^d8a@DY#?R08<\T3DKTM_C<FPNgX3FQ7\VHBXbGB@MN-B
O@bd\d(MUL-W)YN](\8W>4]3@gCQIKBB)19,E^aX@beOYaW?1;LQff-10(0\6FU1
18KR-6(L,bg9^e34E8b;IW-]U-R]MbE7[62B5B:HU+A@LPRU@fd/6edHG;1c&0YZ
5)c[W,6:ac4U>HK<YZcIdK1,3Ee,QK&A2ZJ<#W;R0S,=+LNgLdfZdBL+,bXabFZ/
2#IA)C7]NeWIe7a[H@I/1>U+EM-^Y:KBD?H4_?M3EY?BQ?0I?d^MBg0[)(>g7_XC
L^?Ue)A3S^93TH,_eT((-XPVcf\29P[4+K>EY53E>:f08BWNOU]G<5^c^BJUT#M4
&?c4e<B_?W][PI5a-_PGL0[)7\f7I74V]H7FA&0fF\8JV2C0+aAHOAR&98<&c3,S
#EQL/+NQeTQ2d:E0gFR?/HU0M5bGIa@/T\]5d#P+1=N9,N6Z</M>#_acC)G/-WW0
.,+X,M=ZHF]FCJVReH9/?[S\VUR5dNU]:\+D;e60.=ZKUN+VK&/,0-.1f&B#-PEA
7(#IC2H?@Q3:7>AL@/U/-B,:We.O=b^.Sae7LT+<QDR)8<8WUH2F8\bG;Df#E;FP
VD6.3I#b5^c;A\S#V.+Gg,[ZWa+>\@c/SH;Qf(P9M-):N-I8e12Td4OBO1B-S79(
KV^DQM1.B5N0>LgVYLe)+d3((^:9Bde>PCN.6:))+@+)6DOP5ba\XH]5BgdI4(aS
F^,Qc0WN?b-If^3?]G_eO;;P?WEDM_-LQ=Q=JF8V#SJX0FGBLBA_YRN[\X([:V^Z
_PL5+KYSC7:;[EC=L?VTV7[3=/J\6L8BCBf,R.STVFK-ME07T.4/Z>aZJ_-WVEf1
QQ4^H>)G6_<Z+>g2;[Y>DKg&O1;C3R1g9eT1eGJ1JJG3OI<CHT4K/O#7I;Z+L7[S
?Sf;GO3..d&A6D[&9;#:U1)bI:TCG?02\g:EM?3d[(85;QP]]^Z@1?,MA;,gX;/5
fH.?^cB&_.S48bQ+:Q,F35ZH:;9V(d)9._DeZQ3)/1^_5SXYYGTR09eY@:T1N4A2
0F2O/E^@1b;,K3T;&)#0cH#&[RdA7@)Z)(g#_&gEV^XCL2CB.9@M31:QX,eD4[&Y
d)J<XEB)C)5,]ZB>]_Tc>_X):<,H3;0ZBYO3[5NVQS:PS[cb[<ME:)MXBVG8P9D>
V?bS,XHM5KX.g&G711P;TcW2:=6+IX1-FA)\Z57\P(?.O2D_KH,DV<.[<9:T+fDS
-F8567,.OPbZGC-U(VK8L;bK4@41:;W]^J:#UMTGUEL,DgPN4U[]gIQ[JB1C(L\&
B\b6)\RdBB_P1Y;0N#Z4:EVdaU_I(L?R:O0JC<\aQM;=JR6b7d(S>X<d1;Y_V=b<
AB7X=/8d;+[.4Ecd,=L]f\DHJDBUg8#?)YPW#9+\3YUC_eJdJJ)M5:1?#9DY>^eA
.)T:]/&@<?WYJ>_c4-2FaN]_9-818OI/D9VAUL>8DL4D7RdK=:B?QBbbWcFb&Ugf
DL=LWH-GMCG6_=U=?/_=7Q7SaI>b,?gC)4[&ZR(U_P\<\+>g+f4AV\I>(IgTKR6B
<7H,feMN];YMe&]_>E5J1S9eG8#1g=E)UL>G1=KIYf_E,0(20@AV\;4Z=Xa5I6A)
4.B1gLGB0I,LV0<c]Ca::H-W/Z52ccReI5OXJO8&0<K@>23e@VB/\O-d2Z7MZF:.
3]70JNOUOW9WMFPfgWTP^GT1HJ-)I@J?F8(=bXPX(EHG.?;K\+N2X[C+[cE;gZ(?
RKA67XR?Ma#caD_CLS^dKOCAE:H0@aT\E]UN0X#W-#Y^&S5LFRLgY:4^FJ6OTgHQ
<,Pb@eYL[7Rc@GbdGcW5.(E5+ZcHNDFXg&]LL\.6YPUUHd/RFaF:G#H59U?eI]9]
&3@_/=Pb<;>KWX7^^PP[Sb2e-JSNKDLJ&_&cQ/OBXP.Y>DKWKf1:a\]#M(;5.c>[
.eNIe:e?G]5>?g.C,W?6.Df:7BdP+gReN.WGJ^.2&BA[.&GbA^P_?7f1:BccC8C0
B^WTX8B97]<,><UXZ@4?-294<+ZH3.MdHOG?,Fd0[B)V]0d/M,fB5RE_W#)<CK=U
F>(GJf;N#98#[Ee/FJY13>D]ECgCZJ;FKI1\73a-:#4>E->;<FTeSR[\R=Y1.c4@
J]\f\PbTe08:R+D9IE;11K)P<^?c<;J<f=CW0_2Z+/aXDT\-.^73VD?IZT,3RQ8/
,LD),N3+Y\Q]OJ5/7=a>[<2SbQ1ON0UI)>fBG/D_?AY?Ad-ZPN)6I,71+1)QAZ+9
3>=80N:=[2RG.RW?<O1HN2GN@e.@?JV/&0Nb,J4=\P923f_aCE)>/2^ZTFZMO4:\
ZCG/^X)(_W)RM4/:#2.+B(fX6aF)1U)=Uc\4Q>;2WE=eLB>-)>0G5cE7#)Q87Q[<
.d[#73G02LE2I43VXT00/ADIBZ/a))[FHV,-(S>L0eJM_,>#JW:gQ/N6@OTeJ)?H
FT]d@?Z4]7P^C>4[F)dbW@E=c-WQ7VLQ&P;\]@^=(7U]D;H2dM6FO3RDEZb\NM6Q
>(eY7&Q2;L/E31eK,1WF>dd\;1K_BU=b4b410SIFO9cG@a?>7#8_9/\AS5&Y)4<0
^P;>K-gg-fTXMAeTF4IM@41220R>+bL\>/Mf3T#J8UTT>6DK4S^7dS,,,95MbR6(
=?6B-BR&eU9(Ic-8f_81#A8&EF\CS5:67B2FVQS1QM(7N\E/ECd5DA#PRg<Q^#B,
IF4ed0^>I^gHbb]aaRD73#X-@P&,+OHOARg[QM2[JST.>G,-M^/b0&W_,6DgcK:.
dL(AT[ee+8gDJ\L<\QQ\Fe4Rf?9B#B7V58J8.)4.&D)a^?@-\C2P_BfOE6W=FaB>
N&ZHa\DbG^C,aHMOB1</^GCF2U.,QM[\E2;A]/63I4#=J#]fG:MS4I4OeISVY5>g
UF&?#Q,B?\CO2U2IIN/-@L+@,TU9,,YYDP8N;4[Y.D9PXO[QY?Uc?-EEY3CVODYH
R;-G&1#\^_K,b0f]&<geJP??[F@0a/M6HA:[@-_PYDWL&c_(^YH[_I;S7R4>0MBO
=J@1D=ZUCZK<5\\7.I^M?0C#\B+&-[eK5_(E-M1JEd]>C)EK,Wcb#N4H1^S@@HF6
M01YOY40d\Q<2[C\TY5g/__]82J&;.Cc3UCA<B8;,Q8a3_DT\QX>\H1TOgUML99C
=2X2F(C]c[:-YdM7X-d[R_K\/^^(KY](5d\a9(9g2NGTY5gPL:\=3Z,;D9S1:N(^
-(S6F78[44Y/@SCB4>.7Fdf)[=3(?BR4T/R>K)2Z@1<K1],R49Vg8B6--ZA7J46g
YN+J-aK9T:&&2]NTWRCOTU>Xff/6[]eBa&>1dBRR0+5P\+^:a)_;Q;B:5GPXO:@R
LJ4b8M,U_2]f5f26aV<8DaS9R6/\9\MQ)#W;;VS@W.-=?TO0fe.5.[dBbIR7CO=B
MK4/SAJ4)\_IGbXPO..?2+5g(OVa/KSc6U&<X:TTKg?NU\G6dLJ>N0)gg1E00.UK
W52&^K,bZ>^9e(4?INTaAOEP\aX\3B6QQS0V2Ng1)_Z)O1g(JYZYMXR+6RX)JFZ]
U-+&L9)@5/E19E\#a[7<M&A)K-JJCDBVE2TGKJV56_\##I-YSc?^&b702JR#GEK[
G8..14LX4^QGV,\S-]7F#F^b#ZGD)J#^#E39^JE&;<]NQ#7]d=T(dYCX?A;MF]C[
RF/8HO9&Q;P3Q:3R+.fT6+B0RFcN/g1D-0F&BaO<>C4:UU_C;K.NEZ3[TG(Z?X+Y
]_cLKNa^0R)1[-L.KKb)]>>A[[;:QP>&U:\3YfF8<(Z7@@.gNFB.]D3Aa&43^<b\
Z>;::7R#=L5]dF-#E9bQM<Y,IWe(K]&.>F0<?J,:>B/<dW3[CbZ,NDOdJ>8AcQH^
6[HUK,)Kc6FW6X@V#XgD(8;4N.MORX:4?RD1-6/I0ca)6PK9L\Na84S(ZM]4OCA^
KW+SHdBU=aC0CR2JgXOL4cTffLaD&f@2-dRU2])S7=LI(B5X^_HLHM8af(Ic(g#J
Z@979]f.H08UA>[AIBT?2gPAV?&Se>W0I<G5:B:4Z>g,2YQB[61<C(#LEOGN7?(D
^&=BD(RbG]QXP+>2X7GCZXS2_3&6.,(8K[Z(VLS<gY?CWE&>\+&-EP4ee#0U433;
>1CSJ#GJReJKVX3AP[SCXD+WBUHKT<UM2+b5I9eV:ba#Ygc;1Y\eWbE>Z658d-eg
+H6Wc+EE.Ca>e:[ad(?+]Ra4^+;041Q[T,1XYdaVfMa#^P[SN-72cAG-JM/.P/Te
J_B4@X_Q.MY=dc.QWCPSFZ>+&4Ffb9REKAIf/V-BAUN/\K.?+gP[RQdDdaL\^=V4
A;7ERd;V/ZUDE/W&0H)?]2H-E-0)NNSfPAIb3W@g_f;2EYgQ6<-1g\VFH0ZVb3G1
=FV&:O:SN<RTc/Nc<_)#O-3&AV<)/1YfQ)G9@RE);DaP,?Wg3-&Y@Sff1MVC3:;W
I[2FB&aHeIdBI2V-+W,].=27egU,b[>F-=E<AA]OCbIe;Bb[#Z5J9PP#71WC(Ma7
43ff5B_FS86(gEG^EL7K&XBHVVXdPAZe_=&>LPYS;W_&#6>+3;d5Xc3Z?NGC3QOZ
08HCFLY\:f9Q8&<./Wb<AX9X7/VF7gZ(g/gZX)G:,TN6&H9Wd&Fc7P,@<gTBQ1E+
T-bV2F0=>>L2W1Bg:dGY(LZRF@W\/HEU3OBdgdKM4+<<CQ::_aZTP\Ug?R>+e6Q6
M]0c)U@-BMJJ_W+>#gRLM;COJGdM.]FTZOA,deAS(HA6OLDfBa5CX+&ge:7&0-@c
L@/EMWNX(_/EW45,[/S3]1d]O@b0UV1WDU)\WU.5FPB#X5?:_J0TYG)8#L_BL5=8
g&2a7VfNC@5_;N[[>W=PYTL4N1?HV,d.FdV3HJ,JJQMHHAA0c@\BH.7=V_de@R[,
S(P6Y>9IQ[-FIKD_[IHXBV->HAX98GH+LAA<D9S^D-LVR)5@F0Yc5S=U+>8BZbB4
FR);+JDA:DY(aL_VVeb^IRJc\)NX@FZ(VM_S,3X@+B_5GX+b_d_:RJ&aW:]LgUP_
PDMUVY@(ACMBJ@:F&FeLWbLNg0b/Dc>e6UJIfef(WTbN)Z(=TeQ8V>d=LRdaATg3
B0PUNJ2-2KPE/L1U)fA?XE/(NJQQfJeX=P4=C,>]WN\fALcX/0:RK05N5?DLG4]W
fRXFK]=8+)#I_C]7ZTP<[fW&EU7eIaV1d5^4gH2)bXGbL1035Z+66SI:]#=8YF#H
):81_WFYeGeD0cS]c]O95d]0+>@:JF.W@.=8](IVL5LMBCCeQ-N9>UZIKS8-b;&5
a<93W5,dEK3G:/Q,fY0C-g8.QZ(LKHAHQJV<-Y])4;J=aXR&e<T-Q<bF6RN.AFR5
aSA\@cfD-Jf3bNSTAZE4CbQG&[NG_KXGUIB/V,B4P^1\+/AJ[#8ST\-TW>NW.RaQ
/9(fKa-(>2YZDG8Ba2&GJL_<F7+Ze(,V305PQGW5CP\E]5JXCRK6\NCN:VL[#R:a
;H32T#AB^>LI]dPY53fd\6O@>A?UUb5&=_@DB^>FC4ZQOFOA8A<a+STd^R7]O3R?
DDBPTZ-f<5c7J/a<Ic6C56C-V+>7Ab(JN/<1TL4Uag70?)9bNR=(1ZP3@#;54XUP
d5\BYKNRSb7b)S[+F,feJ-Y@9,IZ#OGZ1>fJ/@a=HfM@X.5FZ.g642N-bB6WQ\JZ
J9O=91C5<5SUQ5YE,_)]6>@ga+#MF\__A&R4E+f(X;IUC5+K+6MbcH=AZ6UXUd>?
D5;C^5Hf7_7H7.ONG2.-EK?gV4E[,H.-.TKE]+OAEg5;97X?UO#aCdd[Y9/A+/b[
DDT2S90d[e1F2-;7C-LYXIFA[GMUfDBUL7PK5E(P_7FE#IP7bSI#ET;9GBH-VcP7
]?1BSQU:^4F:+c;1LbDYWQ7TO?WHF[\,^3gVEO46gg3:Gced&c>2gVP3;I&>Pd+9
75bN1d949=OQDYbcb3B>/W87IG2;6BBE83c[OB[SA:EcSfX94P[d=Wg#X<&ADe[B
gYI>g84,a\cI:b<M+/GJ1Q1HI:O.VL_aVJ7Od)e:Nd2,TL-[73BT9)]JJD#M582g
cf8CMI]^^L<PLN(QUb/^G2dcFCU7NLg4F/-<WMSfA8HL&<XU6fcIS9<X+>-5Y3A+
[X3IZK_eKQWDN+4M<<[P=ZQWLJA<,:0Mag1.4cEPK08f4.2FLCYc4^=-JN6HB_#T
>MeF(dK;@#[4MIg[\\3RSLO],2T\]IC4]BNTTCfgDcd7>)@W]^-BT6:-d0,GK\b(
b3<-]E#DaWYI65N1\aBd<9_HKRCKa]LZdNe?ZegKS3@)?V3JYK=)c[gX#[69C.5(
eW/<E6D7b5F+87+^E\_5@LX&9QDa)3cTM>f(O_P)\Na<&39,>)b>>ReJM]gBa7^f
Na,PW4^1(#LP_X):^BUB9f@VSQ^M<@PS&(3=]4BFHIHfeCWdTQN:aC@H>2,Ge^/Z
P^X,8[:d,>M:KJ1U:;e(]RRA#7@bN8QRY)Q#=c7cTB/gaCGdAL1JeDBba;,FZIKQ
:&B082#fB@.Z=6Q^[Z7.:LAa\f^N=U]ZVI4GMG]OdX?G^&OcBf1SX\YWeVeZ/O0G
MA8UZEV)Bc^.BM,W#dX#>TQZ3D:.9BTX:-V<OAWGE4Z>Qc.2GA.1\#?dLQ\.Q9B;
\9TI+BDP\5+R,ELga:3KT\#0@5/OJBEN(Y7OeP0+OJ]b-ZLK241\bdS#YN;9#<28
I0PV.+#P77^:+(XG_1cR)IYRLBJCILf9d_e7_40B#dPcS]WPYV,V9BAbY86KfX2)
BB,(_T3:bLU/g&3fbL7O492U:0GE+e;@3KeF).XJ&@EW3c,<&C=&0I5Bd<-(3V_>
-cfcS.3_c6<:0d6^:P(_22&0+]_eEN(^\H/Z?-EJS3/a_XN3Ye,G6Sea&B84@[@@
O0.fB9&3IcB+8LC.7[BE+N/>2->SLVXRE(+CK7(dN19S9b6Q=;_V9Q+9NGJ(Z<Rc
aDPabJ.+M_\TK3&aVSaaYRVTfB&D-F.O9TTK[AbSbX+G<USaE3JE^\Q2P?B1G3=,
[2C7/C6.3N_-WdbEHfR4O2+Dc]C+&[S.#1MEg6VaT8:[9b(8OO\I[A/^JPK9#O#5
XbgU,V.X&:_S_U+GJF&H6M#2^cSDSOV&IKM63,I7X0d2:#,\/JfUKS80Z]B/),QC
XH[6M,T\cXR2A/UMbYA\M-)@AD2aGb&B3D^7(W8XE2NL[4eX;Yeg?4a.[L3J4DL;
:&Le4,-^CCPEY=)+=6NY;W6K?0RHG\/NNBJU3?_bP5IfT]eV2P(-Cgc[VP:=[JY^
X2[C5];]8H;15VJL^.T+3K(;Q5I\H<HeA7>(OGC&)+9O-;f<(_6fF:I2@O68;6/I
b5OYPMcT.)O)CFM,+3-b7R:#P-e\E&\[]P(FQWMB=1[1bY\^c8913T@aO7^?Z=c+
\dBJMdcJ46O10X(2=>.UVS:(>?:?86K5Zg&Q(7(+KS&>WC#AJ-).(4/<7C;5/;6C
-\CF&6O7^ZIGQ?(YH[O,>:MeTb3e><^8I[;^5,e4a,f9#AGLC-VeASO5X6c1Z47S
\KaR]S;fL7Y7[;CX7Y,^;LE9>>AN><ef0JaIdHW3YN;YD-5J1EQIJ\9eTMLTB\3g
J&1-cV=JJE(A(CacTg/=4M=VDP9]K]N7N>&fGVH)I>W7H:=b;6<bUBR8V-e1H=8-
b5XLUA]&b&QUM]ZW5RU(D-\_/g0Z4XP2QGNY^1LZK[GJWN<7Ffb=>WYMTfE4ZE/R
WX>N-ITDD&=a<N>1,?#K>&^^[.;>KN:A#[A&JD07=SKVE1XBf4(e6C1&.PZUb#AR
GI:)f4e+EC&/1_(3(_,4B\L&@ICdE6g=EFO.N(SbM(1EN=aMS56gR&)V::b]1]4(
6J&;GdT25\8a;cS)SRPAT#0D^FfVF>DZD9c--@E(:=KHNSG.X]352NVMc44OA;R.
d32a<)c]HV:4)d9OOQeHEN_OPF8.5LX__f5N_\0[<878KUA&X&=;UT5=PNKdJV&V
e4]0AV.5gYSF]1LSg3G-&ZMUB1TC7FG(?SP)-AeQ.?,V;54+KJ\1O\G9WL,T&0H#
^WQ=c3?5V&=f+g/(Kd(+&)Vb<6ZGIDf,VKL\C)Z<&9e2;.K<8NQHeFe6K=]EUAIe
X<NB12PY2MA8#O(WaNB(5CR;Y.K00f-XZG?S@bW>(F)]>EIge[;L,>CH_[J_2H:G
U/T7a?S2D1bE^0)MKIC_V2aQUY#6A@_&MB([)b(Sb/0?PCD(4a]?f]:][UL4=5X/
;J9bE+eRg?c<Y_.\RU-R#bRJ^N=:Y_.JQ@EadA&>L\b?,AQa9.78]#^Zb&W9YP,&
:3VQE:7KP4MTKSI:0.5[8O6dYW:DcG@V9^5KTY9S\GXZ/7##TK0V[961J;\;)(1]
9)W+?dTLGP(7?076b:H7<=-0g4[.,a<1BWJ?2Pe&927aCCEBTcZaBNP-NPc\N;Cf
M<Na7IJ==VN6A6@a#>+@J-GR@F]PSM:RJ933CY&DQL^28]=HEQc3AX\RbH\9^KO_
K)MAb,7=Q^]f_&3NBM+D+0BMQ38?^gG^)N-56VG];#2?gT>/><SV>Ee@#@3)-P4U
eL&@<\L57,)gQRSTYP4XLQgIF:g0>7F0c_=A3C3F#9[4.(faH945F.\:6)&T1+bU
6YNbF87<@aV4#7EL]JGHF7?7PZ./AS@@P9>R0bGR0@3\#1;[RXP#T;HcPBA8ZB[O
+EA@]cYXf/f0IX@1I@)fXgZ\aQ^.cM/a]DVfH)91_8+(A_H^S7c,G69,bC<gO.ed
ZFGc09eS.<BC>,KA+/Z?7ReLb#KX\aX1?J3?@+,Mb7-2&DJY,5.2Q=VN-29GZM,H
F#1OSXFfQB87^6@9LX#B5a:Mg(MT2EL^)1#g#5<NJ[E4<I-PBeR#M\F&Y5433LB)
]SWHA8642-TEFEaQ#33O;D<_2T84W<KV8V,fVaTGgAbafc3fPKg+0;R6+b].3cGc
FQNGCU2-^UP1?2I(>5&fCc\d<TMXgSXB,<18:EV<^G;L9fFX4&OW&;&>?F7S]8G^
B&A)Y\[f;@53UH-?d[N5SR&]H\FaRMIdTOGP]ZYTUg+f,HUU6Qc,3c3,GC.>&D\D
O-CI1(#OPT^+H=a7X0\b2RFcOO:-/2R?;gc^^)Z></g3fKa&<FNMF]>Qc#IN)d/X
<_L4,,M#MgQ:N79.4?)(R)g4B=[B-KW9LAR6LF=G0fgONC9SU6RQ07[)WG\:J88,
S&b\4ZeT+H,_4L=HX)GR0@f0-[ZbLeW<\\#7)O\9)[P2BI@N/5gVEHWI>5YW5W5;
#<Z:<NO4/FS15Z6SfM0O8K3.YEZ+R8]LSeY3SD,VLc)O>(D(fW,AbU<bc_/c-UXG
H<1I?dDgCdCUR;(dEUWMSe/Ofd\NV?6SDZR>_9_g<4-^7SUGA:4UCN]J?f>,IZa9
.\]9ER?<gTN7DaJCd\GB+JB[6Mf4PPC9gLfT,BER5U)62^1J)[59KD8=YPZG2<fB
H(,0F-9]@:M-WaN&-4cW/_0Rc9bC0eZVL:eT8QLFS+cdF:,K[N?CF1]2O8HBXOIX
e9[XL,_:[[JBHa(f#&QGEQ6.&Z+)?TMC\GL6cbNH^NY(.fcR6A5aA.7(#P@aS8BD
^U95IaLOBVg_SP^\OfUUJDZ5VU?L3DH5W9P?ZgVYGKAB:SQ(].5\R-YcN<IXV]64
]dJ1SLAd.Ze9Z0e0+NAV755FA\N;(0_eVR,0-NH>b#4]D]3=KLR\f)\eQfKYAY<(
#<1E[M81S)eF;E/SOP&dH=&S[AB--WHgR>_)HTY^Y(YJ41HTf:<c9eK@H<A&C;gH
BYK27KV1Z1be0eE();4K47K74:E>-W:c3.:<4:PSSB2/YKaWFd<dH9BZ7/644F+Z
3Sd^PP]C+XeF2W@H)+5Y69FA,1@/RES/4f:c1AKe=f\K[G(eWf-)#&:</2SAeLHP
[N9dR3+YbVQ+_>aAZU4OS=.\BOPaTKL?ACK89:8fPI@)55::@^9-5)?f2ebaM][6
C;D@Nf-(2Ed?^8GL2C>d?ZfeP0[9,V<BRZT3@CLHY8_.K?.F&\3Yf/:HLAeO?;V&
N>ZOP[3a5LRP^\KO+/eZYYV9]ea^]=3dNYF6<@Z&USEdG96V1KEagOCCSIc(,L,T
];BZb3UMg928P^(7f>MaI<19=J3/N&S=E0SD&ZR8RT]Q8A\C4Hg.KA+DGDf-\9>W
+(-PZ0b&G3-e>WK6P?5CTV0SN[R>>I.G.-ZY3,EQ\ONY-88OL0Z&P;WaTQaOA[(>
>cB7ARNTX?VFZTR;K<XGB1dHVB+#WX,DPX,dZC7R7=)aa#VEGFVRT9[d]1K.BX_B
-KMZLSJPF7;eB+-4I7C#I[WDJbF@;UdXN^:_RC<ZNN52Jc>b.+b-L8;S9b[?d.B:
ZJ,?:>ISLXRR#Q=[aJWHRIa:bS#]Ga2(NfOB8=A/-/d3P]KO/,)O[Z(B8fU&OU;Z
eVL71J&J2:JM[:C5P3,.LTDKDUYLK;E#ZfQ4AT9[;6d)DK>\:.>U?e;AM6fS,KVQ
Z;QD.NMfA975A-CKLG#Y=NA?ZQ0@<.\TfcN-[VQYHa,JP<B//X>ATCd[eMO(ALJG
KSKYgIU;+KUIX0.>LIJa[MR)7g-Pe^-6^M)g2^c?]PEM+Lbe^bDI5<7[N3A0da+?
J/L]ITS+^AFF(eQC)Ld-W(@U>e]fD48XX6WgQce8;=bSE24e@:N&YXG]PICJ6-U)
:LNJ@UF-09AR-\#G\OUf/#7=C+dJIO^X>4A.2JG#:C@Q@,YB^\>g5;FTXNI(-eQ/
@f=_Y5g37S(C7FJ\EedeC+O8JTf\-[d_OED[3#;1Aa@@<?QdVV>[N@0]O63TA6[e
U1[=^FOAPN8cE-c.LgH+FX:ZY),FT<R3Z3a#9()dc#@;>#,(B>(XI=C/M0>K(Bb=
H4HKY4>5<9?UOV4@bK,^PIOPO__H^IXV6?K]SdJ]OXcQda1L#82\TObOU8d/b2^T
64SIIe-cgV1+?.2/@.-V4QF^a@QfT>.bOcM)6+=e9B9c0C-9.VV0T6<cBf,9eH3g
(TR&=&L&<\0+8MU/#[f.Z2X3.H]I,<WaNQF8T4LWUBcD-JB^e+B3/&<NF,QWfD.6
RSCE6^,2K);MJS5YLW82LSU7fG/TH.9],EO_P,LF)KDS45>G(JTQA,=0<+[dIUg/
NaK7F;U/YEKOgM(Mg:C@KRg.BH+#g4D5>eQQRMSRGIe6+75E_GMPBc83O=:JHJSW
SXLF)-VU1#_S:YK900X4.J^UO1_]5c==)@/VYYMJdR=@XV5ca6&,Qd[2\5-J/EIU
2?W[Ud:6c-eX2^gD@1fFCL.;J__FQZND@[N<.6B#PBDSA]RW&19Gg@1c#1PH,NZ1
5X0)HF90d2=P).&aA^,^b,E-VbC^7LK-N?EL-MPMI(@E[&cQ5;b(VGQFNFZMC^X?
X[K-FD8[9\IfML5MQ9F-d=XH>N)/(]G3Y5;Y&_K_MbY@gRFe3+@eOW0J08P7_89P
)aKOS;S)FS2R+TReL37B/37WH7ET4c,\[W7a.5(E;#JS08bfNAa+D__<U(OZU6O_
/&W1K2L)a=O1EI0=DTJ4_(+_.5.C_WKWPYCCb=^J(-R0<W?<U4c+N9:).#Q6#2Re
6(<>^_)Ha^@G/DWd[.^FH@7:NcL5@E+@9fcfYB@TL#]4UYFEJXO),QF#^.KMC],J
S9JFQEGDD[U)1\3G+9:\(+0@P?9E[B4aS+M?ORRJYZ0aBKf6M9R+)OGLa:C:.Ve>
4[caPTW]:Q(EONZ&9=3Ra)53:+&CA=P_^e9(e=(=+4L+IKS<b&&UgJ?C&?7a1:MG
?ZV5g\YQL/+ZE,9g.Y=<U<Qg=8^](+QW+5M/(8Z\&5K?J2M=g,X2B-KS#Ha&B:E3
0ad)/32Ebd66/Z8cTJJ\#J:K=M;M<>&2E4M_T&89)AX=]/R6;<gE;VR:ROZZ2:-S
QW7<CM.T;;YBcQ[PHd?^0:+Wa9[4a<OWaAa+&+)R\d+b124ELY5^b_QS])&X,G22
UZ^&\>:9SK7a/DfE?=.d:W]P5[,#FUY5<F7K=PfF][gaE-)MNQ0N9f-&3:9d:JE#
T@KMT[N19[:<bWKX^A7-<df\SE(WS;Pa3[7WM3K(A,QQAIOMg=J5EBBNd@7:;Dce
QdP69e4ZLf;7_@fBCSANVP+PZ-&0[@IS34(NJdgVQB+bK_Z<N#/>#aBS+Te3/TWN
E?1JT-Gf]-H(J@>78bUQfI^HQOb0_W.[Z2)TL?T&,G=U21?_2]I>9Y=J6Xd(M_PD
L?E<32ZH_[0S,:SUF@S.gH/H(;PA1E=0GY4&]G#(F0cV?.(SAOO[Sdf5EX79A#(L
L_Y>4D>/?Z,5D/_?f?>4Yg,GCO7[4_1KIM>VV/LQ9:J]fcYdbeB[&/f[-D?XGBb)
PBJ(fQ(8E\/4Q7T3UF5.CH@H]+(Ldg>S3E<,0I^^GaOa3Mbg3K8Q7773_;X2=FR^
TPeAQb/DHGF8a[?16c2/8OP:O,LAFR?@0OMCE81_Q:7HG;M1NH.??P@V=G&>T:a,
9&OY,#M5KP^N0OZJ+]_cV9dWBKc>K\]9b.b@Hg8E4+(WT=@@T]C(T_H,;=0B_U2H
.O1PFVf6QJYQ3D@3&[ABC?;2LBHP@cd-XL5IK1.fK[WOEK&6B&:Z+/X_:+W::#NT
D2Q=WMFN\@IXMYWV/H1<4NH,(YL6H6eQ&Qg55<fUXR#]?6ARf6[G.b1CF9M_-R\1
->]KJYY5dMLbCLRZd7DH]/MLV3Ce]=39Z5N;?<C?.8()22F(@f=YOdJ1,Y_b+.=7
EM/^@T#)AC?RKb/NI_1W-?=N@#W0/XWFRK1>O23.aIQ;>\Zgd[@Y3JJ)3OVBc/U8
Z&e]<cXa_X7e?&f-f^6C7&g\WF87[)#H1,2M_D]M;aVXaW&=U\4S6@N>fSA_Za8I
_MI=<]P=.=.B:10S@>?VP,](=AcaHCCA+)U&DbB]Kd?]g_D9OUQ#+BOba#.[>[+S
B5CWP2-;;0:f7\ZA>(.5Ba.EfNYWe\WJgFQZ#UdH+WCG/gZXK6Ed)_F]EG&T?S,?
[K6)V1M#4UNFJ_J?+([aTg.P-WU-]UVL+B<aEADIIJ#JgO)7WX>ZWAN=@QMI3B.P
BTgG3+6]Q2cN(3Hc41WG.d)CTRJaTIC7Q,]:O&^0:ac+JcI7Z\T;(#4CfCAcT[F/
fQB3K<[M7^7K_E#\=7=EGH.<WfUL)W@P,01PRBRG)(Gc0>DH<e[67_A(PXA)E)Cf
R)gYPG/TX2J/4aV);\M=C7KCKDda(1Yc<LRcHMCR=YM].@0VdY(_5=Z,_Q420b7b
/&BZ4>IcC/&_@,B/6>WfAM>9Mbb\+#[W-\a,ZaM;KSb6\K--#a,YdX2?f3(:G^XR
W?IE]&KUYe=XF9Y&:bQ_P;L-?^6.-)-fY38N4M8G3.H/S_:cZa_E7&:QfTf-BgX4
=]7JSaDT)cIJcC?IGDV\/)9[bSKXN1eEY[d^PEbLSJ9ROBb#(A=Y8G-X)@+<),E6
=:7)J]6De1X;Qf,Ya+(/8gNGI7EO)738V+fPd&8OXUDE5@:L5)-CT61[SHSJ:.A6
.38W+JRDAM:f_8X0[S@)R#IFD/Rg2Ta:<3N#52,K]PISR,eEa-#\U6.)))\3L=PD
4Bf[8G1D3;>N?I?1Kd._F89&8N,T5UU5e(L](#6FV-c2PSV-K=f_M4P@LA)_#(-9
O^ACaW^g-0+QCbTQ5RNQZB(K-+0Pb3b6\PDfA,Xb\X@;e8V<.41_BT2F>eR^NO.U
,(b4TS(#d-53GYG43TZFL51(0S-3D+]ZbH#B\,5<3@LGgPD5T=KR;M/4MUbdFP43
IbN3-1G6,g_8HR.gcW?ACJ^FSQgZ;4eDD/R;B7Y.YS6<@@HIe8G3_bGHZOV+[M0>
ICSfQ\#Z1=^9F+b3If__:\L6&4./<dM#G/aV>@:SK?[;G>>S1(7e;bJN)4?_bZ?D
:cI0N&L<1;KQMH0&fP?fBZN=6b7e?NK,Ka[UJTK,g\I.4dA_XD_>98g]A15c]+K?
N8Jd16^8.EB1\4#)E8GbJT)?Tg=bc#_RMD[,SdAPP?E/KH(905;#B\Ee6+42C_-_
M-PLJZQd5&aQ;2)VG7202U6;L7KNe=.M?2B?ZA158<THS3):D8?LH:BTbTa\&Xe(
DL;3JcH0Qf&930SMN2,gPRRD]_aV8XX9;1W[L0H0E_#Q4,V_E2E48QM@OeP296AN
770cI;,#Y)4LA<F18XJ299S9[T9IM)/91.Rg9,O-E[D-1YB4C_[;DAcJ50D8\\>=
Id&VK]2:8<]B,KN5]3>P.PH_.e)Mb0I&@MO_7)J>IA/P(#3M+XYGXUa[]5e6?;.:
U19D\#ZGHK1eVLf?Q(\e>gPZg.[Z^S]YY9&af)gF1VS?[)3-e8#ab+[#13?ec3O:
D+62CFXfS[/;D](GZg?H9aOT;/IcCAU-=0L.^2L9g;&^/Q8]fFL/I^IVL61TB#&-
75>@R])+E;;PDc+I/.aN34?dD#SUf&B_d3AVD/OBG45)H/g66-IL3R,R&DY7RYPG
@\7X_TWV<:(C;^g^]55D;3_dN<#7PLM,Q<I+\6H-B;;bK9gH2g,0WI5.#BH@OP:E
?P::-+IA&)L/7#7g6BJ6PeYVT6LKeP9?;dI[6.:U.(>aRF9V?Q.AWL5:agN?P;,N
gb2G8=L?OR&LE/GZU]gY,FA@(d[9NFU>/<cC^G9Ucd#LI4]aWX6KRKS&\_FB1gAW
O,+fMNED_:CZ41\QdZV^/N.UI4/g+fU79AFH1eHe?7V0T)=JdfV4U.:S+5,N)Q7G
V\+SC4O&eDD4Z=K/J>/@Z(XcPY+JTEDJU>WXRR4;;T>OGA6afLL<BVd2,W7cJ>G5
@RgI[DB2?G@&PXO@Id<gU=2K\-+@:]0TDN<[7fC0d2T_K.@GJdd#6.f^9+aVI4-U
F+Od\ZS^Q&/#9^[:LC;GUb:\STLgAP:V71,78(VJ-[-EDL2(Le,000@0(aL[TL,G
7T>8>KIb.V,2dbZ8TY:G\2SFeFTe?P/U&+78;6U<fSDKOaEONeN^I=+Ma0B48XAf
YDdgG^L29^,TWEG\.MQNJ;:&bFG^-]Gg)UWHRQ<TS)&W?MIW2F?,7\[F?>P,U&])
;-CSJ3<KQOR_?3g[E[8_\#N#0\e^#)@O:/(@C),cG3=W0UV;9\R/-V9P>WMC9P/0
gb82VVFMd1^L^=F[GAGM9A7IYM.1^=U\1d+0/--H1YQQ\+XH@U&c86Q7+:Y[KdRC
;Rb\0eG110@f,XO3dBDD;P25c5?S^,XCPN:W\77Z(f/D]49YKQ9^Cd,fg^,)9EN,
a7_C3Y-I<MXd?QO3CYX,GeF^ef&a./c&PT/b0Z^.5T,e2+(2g1#T_9HDJHP@>]S@
ZKKWV97U;8\;=<S:560@D=_N]QHRRUBE6]^NIa6bffMCYEIN7:7=69HCQW:b(3IW
ZVd?S6&GKYZABFCUUAF]X>(^f8YVC9^G:LKa1O[HYaZNB?5IWbUENBF1,QcV;L;_
<;d(85D09D(QY]-;,N;HIa;D8L5ZafV1AfD>I[.J-C,;_NffZQSH\YZ(6ca@b9.C
UJK8#.YR_6^@1g/>dZ6.4-(M^5NWBNGP<H6(cPSKWP:S#C5:(<FP@/_D3)eY0:Z1
\7(K)cF0cZgEJ8TKZ-+-I6><Wd5CA-<1F#L@c<?U[E4FQ8(ZGabLMP\84W=?ZM<b
9R6612;??g&]_Xg,.^F0b_>/G9+dKJ6^I)429Ke1=Qc5B7PJ/NA1bSS#eX967T8Q
1d><B)9TAELFO8Cg==4LLGdF\32BQbf/T\C4g:FY0&,IJP#_,N5@Q9f@FXI8DaMB
Lgf\OKK8Zf6cF5/KR2dF&GUK3>(9<D)J1COc_.Ff23(6D^YV+W3FYW?6/7/A:]<(
1f5+2O4fP#MWLXE(@4J_c2F@U6-bGLJSQ&;b<e0\9A[C6Y>K:T2TRB^fgUBaY7SY
L6,5MFXNX115-YAWPBFI\C:YEZT]K6R>;JPU+dUdO1#P3F.M12?,:1J(BSZ>?06:
A1fd#OUHM<4Q@/HB=dZgc.JH_:\8<_OPO5.UU.R4XYXZXYg9B(4M&-:W@bBDW#E4
9U<YcTR=NKJ6#L^FFGFJfScBPSTY8OA24Led8dWZL&K.I<K.H^4FMECC.9QKgI=a
AE\.@@G9FaY57a</bcMW7U>H]J5]2#R7d2_f/5T[d]TP_\8,8S2#MS(@OYcg4YB;
+V3Rg4d6K9&PI^-6,P@X>@(Q\]P[d]/AfZb3,]EaZ98IDQ:>C;f4IKE,g#_Ua>\7
U#]J,)SbN)d\B8.6B)07C]P8+QM0(D68]U;7PJW).5F8(]M1X9,Dc.FI+DJ@;K?+
(MUe2C]X8#/VQEf[eZS-EXJR43f]A@INI5=^2VH<>Ef0/O+XD@OIN.U:.Q/F=666
\f^dMD[2W8a]0a&@2BI+g>0E?J?S<NE7LS\c/:M8a6RXcF@&SROW((.?TS=M0aWO
.7L<J)8<g<f60M=O1;de)>Z>L<[4(CO#(_H;S:;?Sd82d;I1T+S:Ec3GZ87L\S&S
UIQGb=4>HPYMG(4J9HcI+0J](DU09T:E\@4aJ?4aA]=IdN>,FSBW<=(VSCUO.CE)
BPTG6aERI<VOgfV#7@[M]W8S>;KbgV-N5],.2Vg07;L(^Af\)6M:a=)H,)UA)>0C
RfB-9K6_\&bc3Y;]18>=eW+IAPO.>EW?,K3[c7[,Y-VG/#G6g[1ZHE?e94-0ggKD
Pd5fJF9O;00.LDg6H=23=.#80cYWQ[^BO)7D=,O88gN\[GS\^YGEB[JMJ1W&XFN_
cU^RFDQ@JFL#E)8W>]3UEF<a]><0S8#O1A8@QeYd-J@8_b;eKd,PYeF=4,2E(>(.
1[SD<ZP5#Mf6B\TZ?ORDAB>:J[dVS(6@1ZCT0fRW7a0ORJ68gRV;AD]gDIAg/ME9
aCRb,ZJ:,+fU/6V#E/@L]LME?4-+WBLRR]D08@\H>aJ#P>U=b;HIO+GG^0WR\]]K
)H(B/GC1ScNLI@<a;OR;QD-bW5bTSL^Wd&@^FaSgb;1K+@,E[3-#XY4Z[7YL-_8-
#;KZMbB^ZAa7]&MN]_4@6H>L?@&9-E0;LU(_MdB(76cWceO</.3,LOILgK]@5.NU
GaXf92^SJ3DdM+:U@OR1Lc+PFAV8JHI^e]O@,dK1,cee2HJ/-SNDG=.MAV-H5^(9
,<SH_a0CT4EO&X0Ef921H]R/3>R0HA#;@X6C>AbCEff\.537^aK4LX30QfB)W\0\
I6]G8GQ>P[Z12#O,:=Ub;;Qd7MQe]=A<ceZecd=HdF,^IfEW.M:cGD[&W7TN?=<^
-;<#IIBRe-B9)FVDP/VXQ_4^bE+fb9WHLP]9M-IPY8aHTOKQN.;5VR+)4YOSEg-b
:/QgD?ab<8@7#\&_3)]:H.BWOZb+UE9?1Og#RH)29[_.04WFe3:5[5)^FCQHC[:.
J[fT;eJJ5faS>7HYWZ/0)]QBEU>b]&\5/A#0bH>aU(1XJcLb<;@:1L:U=WGS:fV?
S.;XVAMMKd^A/_[,Ne&aC,R_+2W<XFEYf_&^Yc^Y-?MIQZ_5EF@R=DAZT(V@4H5D
QFc1)O:PM79NW6LYN3F/RK,A>^^I?g05C^QK131b2:d;>R_Ad\;Vb/DG,T#(9/Bd
)eDaRg3@D4KM;&>0M8/JWg@DWgJG(1A.IA6+Se4^D8^&gDBARB/Re:7-T<Gf@[U\
dd_D<#5e4b4gFJNJ0^#F5B,_OOCK.CN2d[SY(>\YDA<TMAA[<DK]N6)Z7Ge,>.aT
?WZYb.JgXQ&80:^1-0?;(<[2Le8EQUBcU.B7.aD+c0T83QWOB\)C9^&U824S2;gg
[VX_8Ig0JL]<+cW;?V[=-V)&8g\)]Zd1BQ-;4YOB3b]bC\?8YDW3-K#f)[@,0A_+
SE?^+bbZfW?d>cRR1S97F=9KA6DUXGHS74Y0FU5BRC=2L14,&9+IVNJOJV7MK;,f
N2E31I==-Q37O1FAH6.8MM7?Y@/,/\^RZRc2J0,DDbgTCH-QacC)ecY<LG18(0;V
CS>PTBYJ#\]g:T-;L[-LaIZX0UL([Y1Q&&&.GGIHJ^)H@R1M#&>,^5JSWT^S,9X1
7,[_f.KHH\edVU_/PZ;54K,6QBa5_HO+_9/1=JE49J.D^_R2K.e0d,+HgYDRS_1#
(?T@8YB<\<FTd0[2\M8<;0Q<08.OV@^He/eEI+TVP4>@?]PSf]L[GPcJ88X.Zg>O
1M:c)N-+U>C@_@8I9)_+TO^dF9O\Z:.R<bW[9+JYgO.42,NX1Z(8Z#=:7R;YW^c4
TFNP]QTWD55I?6DN5d0f-9gX,1[D)J7B>d.BN&=-L)cAfI8QVS=-L<K=<1cc;/K-
b.T2Qc;3\^P^P-P.2-#<eD,+Na&XR?WLQD.Ya=,B#AK;V]A-c.R8.JH87>(0_6gJ
HT28AR(3#G?)\=.g7>?0Y8XA-,[^fLY#37D_dW>=KXDa6MAF7TS+:I.N@TRJ4-e-
6>.8^YK&,[b<HfXKT<2.LJM].g\2Y9[F8Se;LFg#JYVIF.V1Rf^_F1eNHUg?.UO<
gOc,EcH=/]X0aGUV17TW2K9/V1GUd>W_PUQ-a:6dJ]U]X&QOV,AR0C),Q<c([S/2
[N^&<_0WTgSW#OaUE,>9M\994-6XNbcQD93=TbFUY5G]Tcd+=P/U.UMD4[VJW#T-
ZaYUf>g@@RBA<BH4P?;gRCFaQMa8ZaR03VPO3XXeU?4.WdQY9a=gNBe6d;1=bJWU
TO[WN08PB6X+D#\C?LY[QQe/RJ-U@B#?cP@X20EV9,\0PT9-):LT)(AER_.P)^N=
9>68Ua1f;6W/LcX&:Y0cf?c_.PMd1f5ZDSe.D/^-BNFRJ)(fKMYZZP0;O[9_=A?E
45(Q\JaDW@;O#P+-+41<@A1C4e@?F37f?CbYOPD]HCMZFNK/:;1LU,dBHM1[B8RA
YTMZZN9cI-Rc]6+b41(=^P,XbGU?FN^gLXDT6Y9AHg8XZgY>O:BR[MV[[NUAbG2&
LDZ26-EJVgVg@7[,dL/gR5;MWNSKbPI:H\H.#_NXg71\R=fVSgPN0QM95+2G2_]L
8IJ4BM8CD)_c:>RPAdJ.OL[KC@,I@YI19=G-eXRBYDc\=6X5.N&_J3T(/H)X-=[E
351>+JFF@3CJ;a\E+K\PQ>3N[A:D?KVH2GH;EgVY97:eLf>V^MDT8N?@K7YK6-S8
1:TITMb9L^aZ^Ba-R]?EDM/efHP20d(BEUZMS-_MB:XYIL_IY4gSU]XJKJWMQ_E-
+0aATH=bC1/]8)+YW/@P]fcX-VE]X@PU6N5>O2;??eX@>Z\LZ^J:dEf1_Wd&-G)V
L31^gaXI3WIaS43OXGJTd;d;AF8577W.S,7EH:aVSB3IC)#(B:0Xc\-?^-R>V&+G
&Oe6YVHdbA0-F40HB/I^#DAG5CI>II=A87_AFYa+Y[DW\>]:FGd&TJ2N+@3e4?,c
JST>RFILEX(:KK/N6TEOcT[NIW,SF\VW1Q=OM-B7#039#5eQ@D+<DCYM2<PGK,[#
U[X,95TD,:.UCFRT78OS1A:IPC)aP3bY0UVRO@ML<ZLa-,R:::W)N)>:59H=](JZ
:9C(gIRAAOgV]1[JEJTcFN@TVf=JBWY<<Y=.a,_B/R^V@J/6g[MTHBgbW(?\)^_N
O+^QN;YQBO1c,>aHf[,7PAgPa9_WYO4F9PR<EP/POceQIJcYD^LXWU<^U=>N=DV1
^+2gG.BWZ>/^:HdcR/;JJ0@8Y.<DfA382@_]FaI.AJ72,_d0\Y2?##UDJ.1A?M1_
&\J+M(UJg,+8X8F3DXMB5A2,b1<2)]ADQ(E2+NPA=Y.8Ce)dKJ-ZTgEU#(]_^.)C
B^S7,OCMW:>4(QNGMR]KQTN,5^9X29+HJbI;5+T/FL.4L#02;3[-.OCLP7OeLS48
4fP)2aKY)TcKMND^I&RX-NcJXU/29Y(3;WZ=[<PN@8JDV_4_2[KVQKFcO7^ATY2e
.@U^c=-0.fXMg=\-VgdTTYM+X:aO1N4RCQK@=^a3D;8@(3a](BL]ec)/VWVFJe2Q
R<\3&=:9EL[K-\O_W3OKLO3RJ(d<b,&f<LDdbX175XM\L&\_(ZGWd4BP)[?B-cNO
;c?X:AY8I=80V8\#2=,7VW4U/cRc.(e.2\5))1X2a>@Ye2=:Y^GILYa)M6Dc]X<:
PcLL7R3gC1Q;6(.>PB?YQ=2+GTTCJB@g;J?=TXH/,J+TPK+7OTUHV;3F?H#fT-,&
)S<#QcWI=f_g47:MN[SW&_P@U<Je&eY2ffW_H5I)NM+0KO7MB0A<;9)MMFE;BbR^
cD6P3:P[:B].-C+(\G5Eb>)8QI1JO(0IC5W-8([Y_X/6gc+SFG4+-X\TNEf\gJ2N
cODP15,:H3ZbZ2.gBE59BCM,ATK)8/U7JPGDJ0N8Y3BTI)HbaX2+f2W>[1.\JN8H
EXgCcT,?7J#IP(_IGOG)dCQ8Z_?1X?Tf[f)2.bf4/:Q0JLQH[/C2J?GWP6\c?_WY
QV&MS7FDZD9SJ[DP8ABV6E1A;cR+UN@gD,6U^c7bcI+QG6:Y@1AWJ<RPN#?ZRN_.
7=D:dFe#CH@W++MIDF>c0E;8(3WZFPHW#c.?V^@[0;L;^,/WJO@Zb)V7I&7U8Q9C
RJBKbMBF-=83/DVS7(4#0U^@;<^N>2cAIN/^9#PRERG,?L@]+N:FLG32A?e5.U#.
\?ADN=a.1&Q&RR1R5@>E2]&3RU[2::H#8I_#M0.UUFB#e3C#DEM6).?1FV,@8H&.
:,9gZ;;^),-U=Cg\,#:Eg=-2b#M[&g)QHQb+&GW(>X#.#]L#^/L>JAF=6:,+FaXW
-,aOTGKYEOH,6-^VOK1L[/9geJ>a0)#9D]:W4H,&Y0SEDFV3^9RL\UBfGE^EQ#@F
^V^6\AV^9=#P2ZA3Z&&<Zf=6<K(>eOE2OEP52eAW\4f:-?PbH[ZW8.;KN;-WM7J2
S\N/,/e:FQGT0BH9L;(V]6Zf.)_^_M--5^CTR#V[0N=Ec09[6@_F0?Y[7MY9d-:)
8X?G=QYG[WbfM:TMT=8:-==T;L#CEXcRc@PRKA4.e5b5;:G;.=>>O>CMcX\3I0@D
58FH]9N-?S><fe:]+;Z:V8>9REA[S27]&IK#7VAc9Qb),^+&LaE,D2&=(g-c\a,[
cAZ<+1?M8&^(L6R0ba0Bag\a6^D,OO\HT;)Z^Ze.1>0aF(gF\&M\5(M#5;J,:#_:
,acGNe)S8UU>5LJN<V.)8,&5U;BK?VcISLaOgPVA[SL\(KH&W>MR5@#-BK@D?7+K
D7-c;c(.TcW4W#YH\QI)MAY3aJV6W\VP1?5K3ZcKOReDXQ]RdT1H<cH;#GJ&)YA8
BLNc<4-3V<cC,B&M^3g4-fH^&3VWJ]E:E6?+Z=:#d3-<0Q\A76R(_f\gg2Oe3-_+
N:A5&X]_-ZQ]4a]X96eQ9aS\N&G(N]cTZ+#JI1=9?I)c^L87:-+MPfR6N6Z?e=43
g3E8M:OG\[M2BQA9ACW;N43O#3dP-2FAgF:g<G#FM7WZ(C=EHG;N-a3Q9-.B@L[P
c^T/+H,=\#6]e5e+]RJa.W;8?=1?bPZC8GME<JL]&+Y,888)?=VZf-UH=6[<LaR2
O?M_>d(AMQ;f.ELTZ6+9D4K54)=8agJT6T.-)g?[ef(5LEb^dWd<OV9a_Y3<M/AA
BF9T]00=AKVU2)2?9Q+/TeZ28A#9_9e8#;Ad7H:(4UD[5.=f-CJScf@P#SbH-[L<
1Ea@X=?S29E4K6GH4b=PWUbN(GD@9LIY#K9,;e1APf9=3]_9Q]-C[]C\Yb=Da>>-
S92_,:K_KAWNSDgA-;YKBMG8EBYBaP&Rb-/JNYgg@_O6O1B3f\/=K^5BO@HRMWgA
(WHUg)]LNM#6X,3eKdc4[-48G&+,,OR\+O,eLRYDLa/bB\K?=4X#4I.&VBa[/Z4N
cB,,/2C?_@Z\aCI?f,UGNN:Z5[]\H9F&49M^_[8eMbE;+KH/)Ggb(c/8,b8:FUH>
?M3)D,Y^U8Fb#OXXfgH^YS8-C:+M<FaE:Ef7A0#E3f#9O=d)>NTKIZJ34VeOQd+G
a#@L]8#(YB-ETDXW>BD+EQ@F(NMW\<D=/SZOe<cg5UL5S+5F@aK0(.gPHFG0+1QH
DX1_#6b-LBH08O78TX0&]b2U,KKHG9O+[V1LFR3E9&8&2O0)=]P],dS8K(?fL0]9
]afTcT024M8OUcV9WfX-U?@7)TZU;TU^8?Y1bCCV/L)HXggN]CU=_\>Cfg[]_\:N
:LK0VYN?E@,b_?EL).-T>[d-1742S[4QSN(.P7?R<(bB9^DTa[<JAGWeKE<?JNBS
HKPg(K=@PZN-OK@eS)XO=6,17EJ=DcSg>MG51G/E_.dW(JK=HKC\e51bd5a[48]@
1-e5,P)a?,&3A+7O5g)cVFCK6[>E7K4/,7M#0(?.BLc9XH-S0WB^,SIfff&Q&Qd#
MR11D,[QK8#7OL;K(8O9=:+<P06@8JK0(-AbJJW]gg]/=&2_VLEM?FRA[;We?^8O
BX.V/HZU7^AXX\gVOJZbO^WaLZ:RMNC=g3Z:S16MECI:?A>(CUT2f^Se\Oe\/bI^
^DLaF]NGfT_D\]OMAU=gZa21d)7-Z9K(RBbNXg8T>21W2b6=>c[D_/4D7D6J;ecJ
&+dRcB8DB6TXAA4F7dHFbK9>#\\dJTI[=g49/N#AL7AX:8H@&\ZM6I]#a&:^>C?&
6VOX:(Cf50[4#:9@4FEPRZ;7PR^9<[+/&E(S9&0PVIaBK45^dW_RaY;12>BT8e&N
06A4USSb:7gLLMB^\+T=.-KK##S<#LDP?C/)#DVZ[9RV=[H9)AE9+1e8\\5JB?L1
/Va;5ac>(5:^?#G@BdM)P]MO<,^X6UOGB/7C5B_R,SIQZ.)&-PB+0^STQ2,?QM73
gM<(Sd_JfRM/KbDB#=SL7:fJT3Fc.N@=]&=7,T)(7-3ccOECY49A?SZ:H6T+19#\
LVPWQ-O4(A-eU^1PT2>ZA5:6^E5<Z@2//@)#6TKLA?)78]4);\-aORHYQOUbcJ82
KN@Q,A,3.Xe_#fa_?dB_c)0e62db\JDKU4:7N&UJL;,-2+LWKJM;Gec=X@M>92(>
_S&]1HEM;X-[YO_LSMgWL0f7Z2WNEYHbH2]\-TAA@WS#IbfO-8]]7M@0BcH#EH;f
^GES&300f@K921;]\JTW&>FI?L:G0RW@B@VAGcbZ681VT&V5YaT6cUS>,>gc5//]
:8AP&#,d]MJ@<[3&_d>>[dI\c:>=M1RJR7^E8?6[)B\2aIZN,+D>MQ&d\J<+T+YL
07C&fOXbc#eBJVQ688#1E.I]Ig7LV3g_#QPKHa&1M(VZ6PS5EYE3^^IUJ<gD<N9<
##6ET5?D?EYD4(\B6&J?7@8S^b,=M-1\F2UD#XX.bf;<Y5Q()+J]A6RPG.29]7PU
Ib)T^;AaK+XGN\g@WWc9=AUJ\1HT0fa0-:(@><37--)77g\ISgE+3BKSH;<_ZBbU
HFIR=fa_5#]>ZOdW0b13WN#?GTUVAX)E>V@Y>D5[)N&,K&N9cI27.f8g]2T=P>ga
5,DUF&MgC61&OU43R<UZ@LGe,BHf/MK[4\R.(XB<6F)=&I;(R6FT,]TM\W>X<.^>
BDN?Tb:.C\GLN6OLL;/66S-:I1BG[9aXAcHgLd:LJ:b=HJgRQ>4A#2F(K#AGU^R[
55NFWL)V>U@=3=71F;/Y9.YKOK#3F<-f>ZVaWg7KFEa1,9AQD5XG6+9fgX^,W2&g
IG?X[9)MFaW/2T,3efZV0--C@fI1Q8&M@&P:?DYBE7Qa@g(XaJ;cJ--a>eXb2[&=
Ff7&1^]5?dbCF@6F:(MQ0(_f<QN:JTZgeCA#T\4I9gJF8_7UJ(_NOSRPE-cZc9Zg
b[I]]?\Cb+HU2[NA9303+6[GVYKTc:#R]0<a//K9MUUeW5#6bOLfY52OMg9JXAIa
]b.Y:<8C.20LQ\[IUJd_S9QAZO\8e2e:4c;91Y0.1ATD^,D0SAWFP]O<1>HTK25)
YK&W02a/8W?7.(,+D/:/9W;]Q\:LbD>PgL3HF>^19B4be_\OG\QM>b#H][U\=[H3
7AVJK#Q@7T\;88e([357OcC_(A?K=1@#/4&/-aC94\H^OZFQKC9P,/J.)T-H^8PJ
^I30#W2+0GbGZ301C=VJG9WN@O>]3HgF9P-Q,>3<Yd:ed2&G<@_@V6AKZK[6B;OU
NK-HLN(T,04<TSaFS+^#ST8;f[?ea9AY><dZ+R]UY7K#YEJ7T\+#-<N43::gF3QM
5_BdS#Tb\A4;6#9/&N,0YB.L5.P5TR;\^#+40KQ4J^c)C/GVD0(:5JR<R2AI>#(G
a+[D;7eE4/+S(a\QgL-4I.F-<:c\<HLU?U8@L(>>X/>COfP./&GP0=+Q9&<6_._Q
[&TM@[DID:gCIOLgV4E<=?\Ga8_,dN\9/@TJ5,(g)B;>>ff4M=Q&/SCRAF+2OcR;
-YF5IRZ/XfdYK1B]+D8)dTO[b5=3WWR7]<5R9PCE@I1T&U\B,6YZ3fR=A^fF<@1Z
Vf3#Z;AMJP7;X?E#-Hc;KT+Dgbb<<OUYdKRW]b>(KWJ038;gC&aMUCPK#7MD6EY+
3(Wa&OC4&QN4Ac\?>PeUKLPJ[?^HbEMEH8#GYfQ5CNFJP>>5fAY]\?U06^)UR(U0
;R)I3D^EW<69_2_HbY98P&;0,PXTO;eR:E42bNB#5F<KL@&H@O^Ze4<M&D4(<ETc
LL3eS:+VHHbUF2>\)6&\41X4?#Y_DMbC&SOS&]9TK\O/XM22:D7+.=g8?a#I4Q<+
(J5MgX.;M3)?0R9#)PI,2f6I3J=eQNb)I8&\6>7N.][VHE;aE4-T<@A,9(+<7?5F
TJ\>A@Y\3LG=]I49K_gSV9#Zea&cO.[8GU]TM&D(9O2Z6]Tc5c5E100\MNE?[g3C
C3QB0>+[Z1g:.A:b9Qdcca5M(O-KYEY]CTO=T-9f:[.2DY:WC1FU5;]S5LUf3?</
[HCeOC&24ORbdJ2#:g23e]3bDQD=?2^:;\:W#&_X27-<>;cR,7cG/\fL7cYg?a7f
&J[#Q0[^,7ELY[#D3>,,b#(_UOGEF+[-(ET)J?80)7]ePXa8=_;83g6,]LJ@f-eW
Ya#=,(&JK\8ag>dTf@?f2-gI\X;;1:Md&<:DN7SY7KRbfSN?DJ013WXH_UGE8KK-
OaGfYNY/OCEGE0d=(0-T9?ed72NE3Y\PDbPBOS<\?d3VaC2Gd\69F/0))^6F0DXZ
A(->CXcSZ^Q.P/KcJNfeH)U#K0U@McGG>3,eWJ<Jb5KRfJUZ\4K8NB46@39eC(M/
GI4HaY=1]U8HgXf&W<UL#d.V<04aRDEcbaGbGGK=<?[WUR[a.edE&<<ZZ0g+F_ET
g@E_<JU<V0<E]g,OY/d=[<We\(JN#\7QCQKf=2B8;M#=eD]_XCIb3B>.3P:0I_5;
E6eYK3I2E@L^<+:S,f09G[;Q5)V-I^UdKgeNU^#g2a/,P(S8XeS3^38fd?0M@\MB
[\:D[:XUaJX\dgC]06ZJP<))b=1,fS)BSE71&ga6)/)SQM7A]XSW71^<\fF01bX,
KNTKMaX;DHQdAE5E=9-]<aWg6=ONb,?Y)\XEVIb:a)RafHgHFf,8K4#-_5]L:W04
f0.9SJN/FM/Y^AEZ:WI[MeCc2D[MEZ_I&Y<c;P5?_[5]3L\f9>>Eg?3+_XM1T6LP
.gI.-6H5R>Ma:e]bU#]/WEeg;(:agZ54;CUC(X.>1?3KQ=WWH6I<^a?RX+LdJ60Q
P:@MQG&5Xa^894eI7I=BZfX3QJ.EcXL/@eRC+fe?Fd+WM:@XUW]PF4BbCM00gM)g
>/9Nf8fWS4T;;4.3a\/.Z3NRLP(0Iae1EF;RBfAIZ-5fAa;8+X7[/#AbAZ-X9IP6
M:1#ceYZA[dQ/3feJWO+[Nf_:KK;Ug^^aEGa8T4^_.f5EQ83<baF;OHSffDQEKNG
9U_4[IX(OXO:aWNI>+3GN/H4Q\fFa=d]HW-=HLT#Y87F;F;(Pd.F@AR7(UCeg@?B
f>B:R(OSRB<=DTEO3BVb\/#1>E,;B4]b/PC=]W/WbJ79488YUFM-09]=R/Y2]Fc1
[g7RQ@1/R;>If#6PZ,^ZP>?VJ6-75_=@+d;eR6W?+8L[/P[5SSQNA)M=g)_AWQcY
4AGd]]>PX33L2WYYMOTT/@^EWYHVM6>gO[<H7ZX;.<ZXWZ&=O;X#936_gF;4HNS9
XB9\>^@,NVMH5C81X-^,:^\TVc)C>=S:B:^IA&g:)gWP;Yg=LMM)7XNcb[P=B71g
.Jf(acd?aXVD3_EGGHS<5@-26<@N\Nd3-dO9NJ(+157<aK>K^;ZgF/cR;0EeT@X3
cCbbX?<\1O>@feNGEOYf/P1I20/a,6ZB\1&DRL\fb>Z(G>R5UgBZUXP\^<Y_H7ZX
e2+1(Q0O44:2J+J/V#^@@a(bBUcb&Bf20Y?T+W6TcV,Q(P\&LKCTAb3TP+=?Nd,Q
92QI:9.Wb<XcFB#;8^^g:#7R84S8ORQY@,(N8LP^G=U@FUHFD^KM5AI;GJ7IdZZF
&[d)eC1[Re=P?=O=/Ua>^E0BF1(]fYCA;,dQGN7SR[RX@f5UID4&K#I-8Y-Z.#L@
=[U[PKMV@e9V/]gJgG&1/V]5I4&@9JFbH2SR,f8/=a?:260b)-<Kcg?L]\@JT5KP
[+38b\Sa2(3S495a+6V9AIDCK##b3EE=9W71SY)XddI9=JCAE1VIVQMYM5)K.A#)
0_=5C-/170>0T^M^I[Q-g<\_5J@1gI#b:/?AReWF-eGGC9fd8bNOZ]_[BV)&[-V7
bN1<XR26_86,6,6;BL[BIKTJg>8AO>[#SN<Wc2(BXCP9+H:&_dffH_^.>NHM@abJ
(8JK:)Y\KNdRCFP.FA&BMS=f^WOJSc\M[WW#MT.;3ABA0]PZ3,4]=9(>gQ.:&>O-
\-CZb:Ja91(b.TNJ@5b4UPH7TMTa?Hg^1cLJUYXMe&TSO/F@c>3?IVF))6_SBKc<
^WH1a=Se6(L+J,)/4L8F\bM.M\ZVE#]VIDVSgT/)R)B+0WR2]fJOT&_4NfeeZTWa
.aY/eRA#I-6M#;5FfObEY8@M7;F/F#[fQA;.3C;A0CNHSI9O7];Mg4Q)QRE91CBU
VA18@&g(AKVfD?[C3LA]-Ef=c#F0FZF+NRB:R9@BSX00.aQNXWD1/#bP?1-6.Y>2
A(NbI2OBZ)Q@gX]NED(1]<5d@/V-a[c^.GW.WM-W89[3NGWgW^,7)7d>KGO0-RML
UJF-@4cD^NZ2UB4e/WE>LJe/6;(f8RgG+6GYU6gO.<W/#/:V+/2L3I81?7e,>UYd
+]#C=Z@.\F?a5bABI2GL-)2JA^>VWNO,fY\=/gcGaYY[=\@V)TQ]<QIUU8_P\O1a
=Y,YC\d+DUEBUD#L&Q.1T:?[K7d^Ub_)1J0:B8I+JDT3[,(O3JEd<F2VA0883JIa
d-U^ZY&[.5VgC\\BbNK)P7C&bVE2@?6NaIbA&&>[7H9MPH_aI/Q\Mb;X#WO6b@OG
:f&P?Ye=d@c(^(FHIaF:VB&4X^:>DC58Z_Y0)^66H5fD>->L&>)^#a+?[ZF(OW<^
].@eC#[f7Q/c.8Xg9T[0?EIZD8)dTPB]cUCHF(WJgd4E5.c),fFKGb9(FL-@T.\f
K3G=7a_ffJb]T;^0&-^-2:7F-CD6CC4PGDfIQ.9J<J13#^IN.7Sf?E@5e4754[@^
Xd79&@2_CHZ&<P&F?\/b0;RB[AW2^HG_):f@&B6&M.[YI\+5C2AGT4A8(\],DP@L
FJ4OQEESN[S8Nc/43Kd&@=.c<0@GU[V@QM-[-QO3(O8)@3#9OQ=[f5bE7?1?S6\V
Ya;?/KM?J:/4D-e/[T]Z1QND4OKM\P;QQ^A_KY\3C293EeR?BJ1Xf6T<]g):8E0Q
4JDW(@Z->RJQII:<Ke1Q<F@N36:P8dPefWaa>NR5aT\L(M.0LV+TT?F=6)D0OX0d
KKBX1_<QW21YZ)T(F_058=XZQ^C@Q=7AA>WdQN>VCGA2g&<EC+&<,3]7XDE2WOF)
/PFBOJ&eYNZ>]JN52R&UfMR067]8-&2Kb1dSgEZ5DIcO.d)CAQY;0aXF<0&4YM62
8F-A83b)@S=Q,36KS-&.X6Jb0fYTFZ^dZ#5+^NCTUH?CX988T40d?ec=@+a(g=Z_
Q]2Gd:d56&@(QFT[FV\5^-MBD2/QHaX_.Z&:Yd<4?C.LSOeGAf>B0NC,02U&V@13
4(7;/C<dCfV:g7SM98L<:GF(.\fK;&(^#;CAdSaY8#bEXRRFGAM_9TfY>:5&eE(;
fdNQ3,ZfK1K@=f=1539P9a=dK34SVY,-+T@7#6Z]B@c4[I8=:WgV],>HUO@2IF6f
\DeC1ZZVVTN02MQ/dAbaHN/)0ff)]^#>P:V4-\,YMMd#:V.IWZK;NCW_4U\,Yd=Q
LH.1DMBTCb1,S/WW2_N?WTS+3eZTIXQ(_H?[_#bXGb7ERQ0KTWeT,I7[34N]IYBU
?LbWbC+C2G,)NY5\N2R/CO1c@6.6c.a.d1>Yf4=O+U94d7QH=JT+8)N]8Ue.57)a
MXUA[#W&FO:H[\NQS[:B)]+O/5J:VfVfOe/-AU#b8.CX^PBDcLc26?f9/I6<<);R
cH?WHJM/:IH>V:^^1G0DU...2G4Cc&BH933F;E=VD:3aIZM]7TADXCb)HZO836L,
J/dLUQ17@0SV86_<7J2QLJHI^D6(J9dUC,b.[_R&9W[))EDBWO/2N0M6A])<LR3f
9cTEMAH6G6<H[41.#=Y6H>_\C)[08EJcPA5DHB3Z\AM-d,d)8OK@0=K5/dgZ_X:U
We9=QJ1(M-ggOQ^GXM0I9F6N;KJNSK60B4A5YE366P/APMS\X&e1:Vb=ZGa8/B^a
b[)N=?-(UYHOBgC7gIWSKGD7\P[Z91S:6]g=g<_9Y=D=;RR4T,UWS,]Nfa->NI8@
N)62eXK3&W/?3NS_WSP7E25,E>VK].Ec8A;4ZVG6QQ,TL-.+d3DLSaSGd#Bc07L6
AVJF<5;/786eK]5g<A[eAOAJ(VK2G_?HfcWgMa<TR#QED.,B@/9CN5=9RP8G:H.&
4Ka.@AU#DaG^f?4<b2fWa\K7ZK6MQ)BR/R^Aa&-T2CP3;<IaCe:K]DbS4WeDB_Le
D@,S+MbAMQ<J#b9ef22bOC:NEHb)&7C&<TMJ533Y&@33O>,HYaHU]HJ#?Z4_=6#)
;+;IeGN\&4S04B/+GH6-=BWg[<73e8E\,,4T56B-8AU707:6MKX9?6^QR2HX<4</
3RKB=c9PTF&3gBK)ERc;#/JNLe)gcaPceMP6@fPPe0-W3C2NdO?NL\AA1)1GgM3=
gEU^:/W:=WRWW^1d-0_e=IE3WL>WL.]2cfUg=,93-IT.9]1,YcQ1C]3cV^JP)[[<
M(8:H#3c>N?dL;#B^A)C-L5Y6SKZEAd\L0GZ+Q/W.P5Z<Y\=?Z_)3KG7[VcTPKf;
c0],<cN&d_H&#?f,a<d2;f8=b2Z[AQ=DP^9Nfba7V7gBYDH-NP@&M0HdLEH4VgUG
QW:_6(34=Mf#(^c\[2^>W@;;>-;DcbU3HKeWP=&=8?/CWJR24SFF>RB>fZH8,+IK
FM6W.4@QH:dJ\-0c\L)J>;>ZWBF+\F;TWP<EH;V=aHabHZ=7T;PSY@JX/>Bg/90c
8aO;YTK>>,f:F1b[=B<gFEMLf>&bc^-SWCc(S(9DIIRe:;,<8@T=,PF5\1:=GJY#
.S1RT4[0+aWg0+<P+Y6gG4DT/J\Ee(^5_2KIASO0/]@H9#WN&-V?W)6^FH<ZfY@(
CHK24W_U01WVS2&RM(.2J2CHf,g)]\K;c^g+b8EA_Y?4@(5-EFIX:d,S1HL25_98
Pb(61PCMfYX0YFGV)U,-^6VND:/1X:XH+T]N#7LU[[]H>M>5MQU\M(S#gP.L]G]P
c&5<H^2VK:R@#QebC5VF:9J43a^3M^?#Lb?F-]ZdOB.^)G5PEB;B9Ug7K#fB@c:U
672DVKMSCWQ;cGXFcT8\O^c_9]T:BIE9.#1G9YaG6Jg21((>e/2F1O8U@M58:BZ<
#:E@0C1ef#cgAba-O+0@&A<XH<^34,a;dB0c&5@[]Q4gS937G-\I:?]+;<^ba=T5
:=UKW,96;,<E5#TXW/0)N3\8,LA.a4e=Z61-;EWN2f]JDR[DD^NK>3)+eWJE^IB\
g7<#BZR>/[>Y)WdG?NZ564T[H\=+FL;NY::OHb1A;/_NIdE4VTY.ET.B54LcXF8[
5YcfNSR@HAUDOZ0:8JMQ12KU>4RX[TIHEM[K+/6.W=.<B9?gZV?72+S20f1Eb86O
aN7[2&VJeDO.T&,DBa/ZGW&?aReG_aPcPM,=<=UeH86#>/<Z,2>[+GAN57MLLF@C
>f5V#NP&F6<3B4_DT.N[]gOU)0H<#-SbR_1>AbR[dMcf8L[gEQ8aG=.H<;Lg2@+H
9=H,6=&33DK2?G>PUMV=>9D,dP4aCbe2?=OB04/3&N7#9XS&ZW&c<?-.]YD1;cI4
B8NA-OFZG.#c#)+\SFLLX[EA#CaH1-O)DV(.P0cP>@<=VLd3L+VH<6#2D-JdR)W]
Ke(6WAJS8R/EVPP-[^LHVTaA)P:&+1M:58f)Q\Q]VX^gT@gK:B;]NgB<L,#T5Q_E
]2KUW0[<N5ADf79JeKaXI.5>DeOcb@Tff^/e]XAB\1L=0L8\F;38EI=2dYR(@dG2
BJC@R3J51/:EJ0f>60&\Jf.VJSPf;WR<KMb3d\@4J>1U-5_@d<8Y0<7P4[\4V/g?
5^M&1b;gaW6T9ZBOd4J6HI_[-PV&K-+^ZR2@aS:X:VP9FX9e7,V=ITX2JWg,/4]6
e;)TAIT(<^,N3>E.EW^f1<YH5X0:RbaG?MGI/##Vg)b.^C\\WX<\K2YMYP<Uf.Y^
[CW[5;7]23a;7W23R)cYd<]3fV_Y+-99O(b+.ZZF/CL(>K=bBXO6:V]YZd:T&C29
VF3@DbQU&?Q=&+0d>?1V/Q/0ERGN-R_-2_/@7Y/BKC-\Z.OgF4Z2fSFbaeOJ1gK6
)CICZ<IK9>SW@VA)M\^^.N0X@8Tca<@gd#XNd<R>(D]O>;-TJ4Z\8:Y1-[XT5LP=
RFUGIcO1G65T-C4ZGOCGGWP_#cG/a[<V,^#A_Ue2R?+Se::QF2^-/VfPZH\IbI6U
d.41B+>663<(ZN;]DD6WG@>78LOM85,9?)\.>9T4^,gMF:P?X2@MS4S19dNQfR@J
V97(aGBM3HIP]9D;a5@V#X5RJRd@&OXMIB7B2f4S<6bTG\dP.Z1daLR./3eUb:.;
+-HQJL935<V0CCbFfW1fdVJ7]2@^^e3]-USM-5VI]aLJ98C7T@,:KbWZb:VNB^^\
aOe,b]1A9&+N)&9Ge9>[,:g#@B\>Nad^O3-IcHZ[B4D<)YGbX?J.;7d>f?19Q^6H
OcU]RR74I1JRG5](NE-U?8R]WD>GX:=\;E;2L;&S90.^U4KQa/C<92RJQHLU0<-G
8SN+7X26dGT#beUc_&<?\#OL1H#UGf+W;MO&8YRgD>(3[(H+:gR<gX(WZ+Fe#76,
N>^95-VcDR/92=P5ZeFf_:.Ma2B08/OLd[WAe.MV2\2VC&-/J&K0ZGGa4&=?f;dE
HFMQbWd#H2f8FN9RUeW)e3HJDVSHFMMM9\EaNXK=R:g7CbA=3F.?9d_GAWR+.@Vg
BK7M)UJd8G]:)475HY(<]#A<baK3AHdOcEFJ5HCe))<e()K(9D/fHKJSS@)U;W[O
AEPd4:6N2(f.aOeM/.\Y?6+.eD^T&@J\c7Y^G?H#Cad#[O>X;G>YRC1A5fF_eb)J
OK&Zb<ZFO1RY:T=_>SALN;WK?)5)De(]W3C\c<M^P,LL,5N2_S/C@#@ABgO+YYAS
#?/DgF<.0M32d<;)JaC>F-=/,41gIV^Hg9U/@_)-AR_AJcDG_FJQ/9#>X5Jc]:5C
Bf)+5Pd.aU;VYVA>E=OLC?d&J\9O3a,EaAgXGZW2YR[c5W/0c43fCFR.&bZ-TQ#[
e+b;?;ZM;,#HJ[\;EO,g0L<MN?W^RN3ebW#;ZeVXQ4W<RRHDBb._\Z<#6;MdUN-N
JL)LS<ge@UJS?AIRNPZ@d1T=gW)dO<gX;<FZbTc+:)J9cdYDO;Z:BV2_WFbZegAB
NgML,?Y;ICUJXL82aC:4-^g:2bIE/WXVTJ)T>GQR9Gb:K1JS093@?:.&HRI7VOHS
[ME=0cZ35<b&8K-^IXGdTW#5=&=G0NN,K&6VOSS<>b#B]=b;[2bN-XP\V[\,e@W[
ad^CcS&;\gJ=-R.E,?:Yc^cC8YH;D0,]46HSO.Ge1,CL\KV9,0?PAQ:?7]1LN#?,
d,JD037<2=((aYcebUTgNcFdHL8&PWS+)ZJWAR&c4YbcLSH,#20L/#ac8N.2_aVf
f?_I\),0N#OTN>EWWVYYJba84<GFRSC(3=G^NHHeE;M^,:3X^&/3/6&c#aY68N3F
/?JS@Z5-b[=Y^@.-g/?TQ#XA+(SfdBNBLQ)O:+,7Ob8+;^g1=Y+SHcS?XW)dSQ&7
4#&SM<TF@H3(=^fR6;OW6A:^)&W3H)@8XDLS5=V9Gd,CRW<UR6ag3S.Q\/Pd(>TY
3g^_L8TI_^CB]bJD>NYfGSTJ-P^U[Ig?BWg)MNA6g2KI\[SeSaF7]W04>K&R:5]b
1FGg/,OEaK1#&2Y5)WX5OdcVKO(8TcOBH2U#-(&9J3<9+Q.YQ5f(g:(<Q9aZf756
N_XV]QfW...M(22b&P&Ya[?[?C>>)=FMUQ(d9R2OWKMHW79N()(.Xc7WN.08;HXB
J,W.J5cUEE^K\Q&bDVR)Ne2S<YIK8JPaQJG]>>F&-O(2U^K(J7FD@8V,O5L@aW@<
5MZQ50WMb[E5CWJZd.c,L#)5)&YOSJ^.RM_KY/cSSKff#9^:f7<Ba5[Tg\Q]Y3US
L@U[T2MNZK;JR4d)3<(1bE?BGKJGQX1:K/J10Ed>>UA1M?-T04eF3ORV<.S[f\I1
0T;32dc1WV,JV:6Q]2A0<K()WK]f3-.3+LXIRVN3&6G[F:^(c+G[)6H6\^^b:ARg
+AI^4Q?0T-e-#364U5#(K=LKWN22cfEY#M5=-TTMX(3&.M\J2fT6DL^_&aQHGT21
&4M#T@[&UAKS+Ge7d#->YA]],>(WVRP7R[&J,=GVD),Z,(Z2V2N2cfgO7^G5?Z0E
c&4F-AK7#A4T@;Z_ARgUd#DOV[;QHSGB=#0L./d2aHcaY8?.VAR#1Q1+Fg8P@_C6
.Jd\E9\FY@<[ag[GVG8>;631fcgN)ID=XW_H6BM[fF52e&74_bE#dP]SS_?R[I]J
XU0;d[@gb+bRG03[83JLIJ2Z]<\_(FSM0),CH7UQ;HS^;6<CDgCVWC\M-V4(FK(_
5-bg<<XK_4,QI3M&AKCdBR.U[K]/?c7PI]=K@e?=MK)2,aL[@1c+TTQ.I:d49QXH
U2X)>[=#7</#TNAG@QU<.B#,25)5?G09KE;P0X^fQO7U9=fFdH&NJBK,B#2IXB@^
dH23F6W?E7a7(]G?b[cbN?7f8^MF&:Oe9O2DA]2C=YFe_Q+18HF<8ZYYZ)W8.XL,
6R28G+K==8@Q0.=6TO5cId70R=5#[.R3CdeWNZE;KJY_V-V5_-JfJCB3;+7BOCa+
#,3TEZ/35-<P,@Nd;+W2X8AAT_/-D<SJ;91(I=Hd.VX;G#93J\34CFFZ/UG[;XU&
J9]WO+3Y/P;XIIaLBCFaG^c#4P.cC<1.[)a8392-MOOI:]X\6.6Q>]dge<&/gb?-
DY@gEPbW5N</)SFG>+/b@J\6KfEe<aTJ(1F(2SPQF;1A2Id?O^PM?+W;-\1gK?I<
&c#Q0(7IDCY(U#H-If.YTR_2]Rg6F_JTbFf(SF&a-IOV5K8b<=K_/\+N@>=+W.=0
fb5.HH@#V5M^D6U;.#dNV<)0=9EFc4e28G/3-G(PW5_DNVa9Z7P1[6FJc-.)IDGJ
0JPX2MeV1D;e2Y?(TNVT85dYecBd#L?]79\Q0:^4E^#XA3>:91eUTL:Ue&0#F,BX
E^SI6[fAV<B5D9Q:6BJ=_VVdGR2AF()63gfG@fX::E)/0TRH/G(&Ka^JNd)g6I>)
7.A5C.J1].BU<RgbKM?N#L/K8HY-OaBC+b(I3X@T>53.Rf/(NaGMEcBL7,LD4>-+
W>]a4+#OgO4cJ7_\aG#RPfBRAPIJVd(-);V>2ad0EaF<=B@1U\;\99BPETU-C,b.
1\69T2?//REbFZ=AZEE3=K/Dda#(a4@C>N>[7H#M@1:21,5Ne^S(J_M5BNL35CQ8
MYY2@3-dcQKQL=abMb@1g;D/JEBC=5;H6[RD>3=RI4D:@VG^:(4FQJLMV1LUFQN<
O0]L00F\39cKJ&-5]1.5(5VE7JWKMX8L#<,:O<)A1a\A5M?PM6P8(Y]__WWcV&&T
K(XcG3R]>eMODL9dZe7f+.)fD]fT,aQT5A<X7C(aQ+RW8dK>(><\g120I?TSC.I?
4D<<[c4NY<CJ:96\W6KY&R]&YUB9,+gX-I]J_#4Ub=I03d;>e9V6RBK#^10HLeM#
NV5Y^fRN&TTU;:HV4^7>fTPe=UIN/2<&KfI^X#ND9XWW?YS.WAeI5OBN&8Q&QWEK
T4);fA54eGIR4CW/VR=e8X?CW/[EH:;5,J#>-Z_a)HNX:UCWN0OA_A&FUIbZS7(-
-P-,HG+:3U:9)NW=3a+g7_cFYG\ZP)b:e4<:_(X=+Z6#W_bU8Oe1(EGK^43^DJ@B
I:+?8^IgN,(d1(Y)eVX&cfeO,L>6XVUJN8-fcQ8NDSHd,O\aZbbYU8D#GS?/ZSc^
@ZQ>@U#&]G7IDPU)=G&B&P:X4,H+1KSHXc,RQaXL6B&>(5P+C;)9/1_7XV#P/ZE3
c0GQ7-@VSaO+[g\N:CN8G(RT[DB/K7MB]/eEL?92,R\)6MTF>.>2f>@7cWSQ&[1/
f9eA@D7XQd[;fg7e9Q9a1fDM2bT0fI[I4>MK([Q.]J8@eW,6?&e23cKB:8X+I3G,
=6[[>,+F)fPR.=>8I#H1>T<8[gGgB:Pd@,\3JONR4167U@ELcHE<SG,TZfce69YK
Vc\Q7MgG+Y[,,WV2MdLL.+d[BK(IIP)LM0-AX3\CH>.Q.6Gbg#@[cU&+[c76WI:9
2H20^4W>1Y?EJAeA//S_@f[0^VJWH/:TCe]EM_YQHGb(^BJ@U6OZd@,DcB>=R^]1
0X34d1R5FKc6[DSFQ&Kg[0_aZeRbCCT1+@7d8QggP<H5>]HQf1#;=\[I3:FeM4>=
)/-KI953BB1<4D3/KY&<N1)7E,4W9Y;;)D:@+W\a[DCaN2YA?^DFS2cFDAWOee(X
#.2.@da>gZdb?>.SY587EGSa?W-(N]-K&F&7B0bW0e/V8bO,36TD;SY:_&Wf3VU\
L=MSY]^0f@GBEQ4/T.T.b^5Y#52=C7+YG^Y8#K-:eCP=Be3)S+FK-eFa3dN,>)_K
SM(O&)X7]3]>e4ONH2GW(03c301P>+CPRC6-YS-UW6,e<Db\2K6?(AZ@J[NHQ53_
QFfc(XFYQ8(Sf7,#]:<X2T=KC[1Yc2OE5Y0,Ng;a?^WPB36D:CZ:6aU]c^_Ac.V9
1gJMN2\,8;fP<S?4B8CWOAOUN3)4)S5UWg/GDMXAAI79;/df894CG8De,C1db<-=
7Z/]/_YU_\XYTOHG7B3ED<;C=^JD^J-W^,[A;<VZ?QE0V_:7_MG5,,2<CgXYF,7X
NQP<9T#L>Y?)NT2\;eA0^W+Y=B;G^IbaQ,)57@D.(T6<[4RMS9=Q;H&1]T/4RD+7
UA-N[c51[=FMH?G;^;\T)-,L:-8GHV]f0QfU@EH]WX-_#RW./@bZg-0STB>I+BGT
M(aWDC081H2O]+e[6=-YIfgf-3fF-T.8;cCEbb6^N6DgW]9_J64V?Gf,DE^b.?UT
EY7J79<P_WaEL6.[2IEE@ZB:>T#+=8+4IFDSd=fW87#SN?4a-Y\fO[?D&3M,_)0V
1A^T&4+NL7/37-CO_(=\&^NB^XecfX9A89F]7VC:J:PWC8/e3EGD<U5C;E2fXgX2
DI?8.TMUc3+YOeSOd9(=[A]F]4,N:/U9CVWCA0F4.^U_UM5bGULF3FBaQOX46XUa
,G-@aN7]+ZMLSY2^Y-HWb;A7V&N/Afa\&A_7Vbg_[\(c1#P=L33_Qg/<SZZ39#Ig
fD:QD,Ne)QTIN1FLfW_H27O2TEEEEME_I?^[,_O6IBP8[D#R#,B@#XD2B;(ZH9KS
__Y^?a;I1f6J2D[T<G,cU(T2H:DeOB,b3b.GE,L(32LT9#C46NaNZYaIMX3LXOU9
Xg([E_S7@7[OM65(@[9HV_L<Q2KJ:=V(D]^<BTc=gbUJ3aeLg.S\,\+ge[/JL8_7
eX5+F,87a>9#]#RFR3Jdgc,0.+,O1UDH^>9?M7g-SdB:gQRQQIAaBc[ef_9N-?c_
]IVg,Y=0C8QZ&UU6Cd:NA]f7]3Q(PE\WDaVN52e^J6022P<1gd//Dfb8BSRS6QV;
Z:_G6(>/&LdCHT?]M]DSLf6K]2R;ZX-[dC=ZX0[eMMZ8B]LIZ<DfV5gHA<;OaEDC
O-3IYQ)(-3=]7::HBKL^1e_J]([H,5&f.=#EX]_PJUZOGfQDYA-QNSf<MJL97E#?
I8dDa8>NC,JO:bS/&4?e07VWcMT0b#:(CYY&T6C80?[Cd3/]Z<5-ANP4()Y2@.E[
fPCf30:fX(9L.Xc>dQ=:cU1a-D)[VYd3gefX+8<dC-E)/;OG893P8KAe&G-fK>+3
J9SID<.VJ-PQB^(a(1+W3#?]9<-KR7XUfL/3K>Ia:-Pfa?:=,51>)8EE3,)<ZdT-
DS35,POZOTdfZJ;2]^UF;?bZ3F-H7Ga=BD)8?Jg[WRTDadL(E/:O/&+WK@VM9CG,
H8,265+1+5]29&C>f5>b5LZ/AJR(a8d][b;G7(VIV.9DQ(QSg:+-M@(9:N#G/NfP
Pg]P@S+8Q&5^09/5/7a:+6gZAJ5<GS;]57^8fO-]1#4e#a7/f)R21-aDQV&0?X#\
MG:IPR/7QHcg9;c6)0LTUd^D,ORBPL.QHb(IYV4(TTN8/WfWQ-cOQ&SK,>QL)e<T
:1-O?-9gZTXMM&\Q=GQ9=17E+)TN0c?\2gSe6UK2Ueb#A;2L7[D9cQ&KAL0GCL(?
g40I4ZRO)9Y@B@Q?Xa?:ONcD(9P/e5#5LK6-I:AaHe)9SZ0=I9/L4L5,(8F._W[2
0\)WQ4aFI/J[CC-Yd].CUK:#,D<Ja9+@<6dc#HFd/,;SB0;^A+:\P2a,=9<NAQeO
Ib>,Sad7WOR?.5aBV3X9&Z&&S^L)+56IfVR21#S:d5.a4GY].6gXPdcK):U0(F@V
]B?HBTYWf5JH:?c;[O8b:AT4GU@5)U,NNSE]V7ZVfQbPVcEOH(].N:H</0#F)Y05
\UgUFgbY#V@6>cR4V,^,M>)B\>4W:eeY\2O8CEE/2^2(396WA/:QX29QfdHP.<0,
OLfCB;_A+g.E(Nc.;4V:FH;JIWe^[.\>2E)#dg0C+[4Ng01)T:,X@4TGI4F(+HMb
Ha#L___c5M5a#]BPKA1Y,U6D\Y&eN^2E9H3N@c>Q#aG0T7&YGX\c1()Id)ZI/F0?
)2BM6S[=#Z-F9DKV<FJf,QGe=+R(XfM;.MfMOJ+@25U+9,b)-?X]\=D]bQ_NE4&H
?Zf[1LcV??_9YeLc&?JGT9L.VL[@>S6/b3X+)[SaJ_;A1,FWBG_TC1c)A6NBf?^K
-K/ZOUd=0Y)#dYfVV7=L#62E)Z,#^0fd[Z\-?aUg;#;PL,P80JDVN<<:/\@]X?F#
@/&5YCV?[L>_+H0UB7V2TQQZ]_6cLU\<0Dg5QGTcd)d\X(IRb4K7+R(#5bV6g.#>
cIWG,1Y]L=:E.[\WBQ4DS?SCd28<(OgLADIQc4.PBYG8P:=UK<N0<V(d28W7e^?A
-36)+bGKFV&KeHR10A.>E1&PIFB(C&+Ya+Hg;XNB[2aN7]fN;)\T5SPFAdB+P)4A
:CR\d@)@KL(,KWT4J>.9<ga]1S/9:GWMOgJFFJ4,6NIOPdW:0=<G3=&:OHEGENe3
ZfW::Cbe,b\E5:g]NT8B8MNDTA?<-42=c;WAC)Gdf+g=297-.MK[]_;H>E8D;bD-
B0OGQUJZX<I,/K[<6&>1.Dff=8H?TY4b;fPAeGW_))BXHa@SFT>e,99OBNYCJ/)?
^1JVBH;7@d7_/9fcO\^d4P.gQ9UPbIJLcQ?ceHa.cWeMKOLgI#G;2)F-:KU/I?FG
@NJ]7EcVCeQY)JGSgO7)1UH_EXc&.GMBS<S)DJAFY.2SYgZ?KU2cTMC2#C)V-C6A
PATK\BG4;\4:??GA+?-B3V_#A[?SMJ=-W@e]OV]B)KA^;3W(K+JZZaf78L431+a[
N\E6:/Y+_F5I7d#G]_U22XK1/URNK?:XdYNBQGa?@ga+V/f+M;0.4<)WPM<g04]_
Q&7S^G1U5S6&-T.S)&3^J18S#(@I9Jd/#+>T)(4.baDT#Z9HcSL[[PZ_0ccd)<W_
<5IEA<.4ZDF_LF)8RS&_)5<25^DKId.Q>K8>Afg^C?>)E04_#bf=IRSPS[]3.@e>
IGNYCL?NeW[79+R,b@B2LK0PGN@]963Tg9gcXO]1eRFGNGNZ8&TYA,[,G6.3(e@1
bHMY)-\V2<)YD5NYcW/[#8)4G8=>?Z;MY+]>6aA,cTL/J>Z7+81cG;]]3JLTZd6P
;>4IM?.PP+4[gC(]A[++(VKNC7_&GU1F6A@;9,1W2-A5?9R&2@AQOS\6>F8M9H@@
O_@7G&2ZL>/([f-R+RIO2_\A#fD0Z:;<\6P=#dK;RJ]MDM=:c&J^^FT.?\S=_fX7
4]P0:I6ZFg7>VG3T@(a9AI/RX>@;QIM&3GB<e;5@S:V;,f^[,LG17I8e&J;?M2.a
N35NP3Y4g][/]->1dF\1ZP@8&/[]Ff-#&K(85UX(;HcXMS)]:ZYeI4AG5]TU.X[C
T0V:?H&+CZ#(A<K^:_XF^\Z)JdR^Ze3@0U7/U^Cf12;3?6JJ1J<B.RGE4Ua-&?=G
Sc86U&U=OE,8ZI4+V9-Y=#d1SZAJJ7IH;#7U([HI[BCd_d8bXI17^0[97#Ngd]OH
7:K0O3OV#=1SC@>/=):G:7->_61eN>@.;Aa)+FOcD9]Q=NDH/)#^7Z>-SJWUWL=c
U\:bFDbYP>CT@)_D53=^41M>&^8_[=]KN:L910\XX=:QF<H&RN8X3(@263bU#U83
+L?KV:;de,Qb,Ue4#;R#1DD>C:)?\B=AFN[]9JH,3S\I+/9CdY6;4&dWKYW2_&:@
/5^c6AX1?fPNK1UV?B(PRVgfB4&Sg9U#0RA8#MKGa\Nb)L>5WH23=\@RU(c-M,O/
A(;I1CDEZ:#QHZ,1;e]D;8,]b929,D/VE).]E(c)<]+T4?FOfbZSWAE5UW]1e-2d
0#:A^0J>7cC6K==PS^UX(^A_^,N:Ac\V9@6[^M97^/?>I#.gI5MON&;+B?&+_W-Q
#POg2=+MB+,ZMGcC;=&RHa(R7PH0XDUQ=OfTG]XOG+VE:V?AH_A,[_W7&909@P5f
;T]GZD5H-RLYb5X)<8#0B#)/^R/F/;<,R=9e232CSd@/8\c<6OSaJ,KRI=8fb4IM
R>:EGHVBYVI)1,0K.URYH20.]Je7=BfY3eJQ^TU]@02;YCYZ58D@SLJ,CQF5eBO1
2O9S,AI;S>]M7^M,VV_P6Zg)>WRDJ9J_fO#gVLGY(MgAa?a;B0U^W77+M?7\b,N0
a5?dc85gOOKUbUR>69,XdAKG_f;f(G:W_;+0+=c[H?GP<:7H\:REY(5+fX)Yc&cQ
?_@7^g<_XY\U5_L;(0+A-g@\aCNNL@4S[Z96cGN[,ZO5\XaH6HV\UM1&1E&D9,0O
IMA5&?J4f29KV0(PM=HQ9QI^#?^TGMS1d^;[aaZ]&NV+JIA<#Z]CUX\R75GN@1>c
?W7_OA/P6f&3H6E3BSJ1,REV7X@,#a,_ZHg([fDMOPXE7eBf1c^4CWS550,fd17=
0^M^^@PGL[APR^ME-B8Eg:[Z(@4Ob.dW,)CaRe-L6/W6L.9+3YZbH+TG329[,83]
JAJNNF\CV@c3#dT5E=4_O4,D,+9-BA6g78>(VP,3\HH_-<e3EE43e-&5I8@FO/bJ
I.LNAGe[)(9FafN5f3PWT76+9Zc+a.[9XX#CbK0#Ee9CLdC)=\>CZ2#/\/72/W4Y
\&XZUgT?8.IZFCMf@AV7L56O]fH?4d7V&J+#aXC/>U=+8-YS(=9Gc[<H_#+.#aI;
#Y+B-5gFL4b4?</+dPHVb>[SUK;M5Uce13Q/9Of&[Tf38bF,?X[c._1&;\ZO9adV
6M<BF>S?aW=5=6GJ5#^L>(XU1O^0f](@bX5SGY_IGVQ7fHSD3=(/9]MOCZT<?36(
_P,/?-c-F>X07-B]VE+JH>PF#KY;2<QWH-.<K/9WTS_B:&B#_8.HgNSag&FG22=L
)3S9\,a<JKf\TA-dTWJT\D_5,]X672WXP<9\YdUYCB34/+H_?UDSM8YPKHaOd<XY
=?L-7.F+gNH0f7Gf>b#G]+(Z9U@dXJ/C(T4.)GQG5KT3#7cf;\_VW<d][/=_+-g4
H>bN:(:BcQU)=D<0B-B^I;f,DO@;FI:++g&Ya1Y:KV&6S1GA@gC.?I3OdD7/;WBA
P:HU(83W.0HED6X7d2HOTL3P-Ca>Fb^0T(7OS@7__=E0@EZT3-1)N5A0ZWS9NXCX
U(B1Ze6ef548eIa/ITR_D)38OYBJ/M1T6b/F0IcEJ,DJRRd918>GI[cbfDGNaFZ+
^<]_M73[2F[ggSSaZZb_]/_F+S1ZLH:Z(CM[4d_+b?WF#2)XZ\I0CK5Fc^62)DfB
g0Wa)D=c3gR@OJT5f9KgG;(24EbKB(_(JLT7@.YHNCN=>]/R(@63M,:RN.eMe/_C
66?cc=MSCMcVG7@#RRb>bAW/975W9@9G9M<JU<96[:U=&#Ee]&:-WVYOS-P2\G)Y
HTS4XdGb>ZR)HY81TDTgGa0B6F3gL9/BcdbTSWaG:R?J\.0GM4G9cEbb(#[Y68GT
5,Nd&+A;8db]cP-c73+NM)bR7e6g;HA>SSM^VB[@.;JG,H_K5_:J?b>FI6-;.ICE
EM.PAQU@2MSa)9e+R2KeJ)I6#1Qf[4C0>V@,3bGDA>(9J<V0I/Sd1E]G=VfV86H=
WcbYQ4(&2>K6(6QYKd^UE)R8(9KG6dA&JH8A]0U-,9WLb@#BVA5P:M7=(JQ+EB]R
H#dVEI]H1X0g&851R;/T)aOK10\G7<b@>@IXT7e9b1,VJ+)?H@gXV6;fb0#2SVY0
A^]8U-eW:UQIJ:9eW,H\fa:[9CJ^U6c<Y+]WT84I]H)R2d+8IM8>LL3@D(=e0CY7
7>X3UCJ.#V(K]N@RS?9<]=64a@[8PbRObWcbU5WaH;?Y)ZCL8_Z=1@NDX24)]1T2
ddWc+CC.6baG]?IbHGF:AQdcQF[M_A7XOgJ:d,HF=6:C&&ZQ5U\[HU[c)dDgZ+YV
R<.WA.JV[5F>U+BV3&_6+8cMGaWKI7f6ERI_-G\GagC8:7-M\(GNS1)Q@,GZ\8;d
U6VROIUTVFLXb6Ka(I-dN_0@K+d&M2?^QGXK5cN,:)S@2?@.fd@>@ELZUG2K4/\>
g6V&W7)X4_dAa[/Q_JDd_V4MIcRa])f;B93Z[d&I:a@cBR(Hd4F:NY?ZDfL?KbA2
5ge/VO)#<b.L4+LZe=cb0+=LAUK8^dVVBXEI4UQ=E#>7QPf#F_UB>(/_Q8b-g5]a
])O5E(FL5Q_L\8YI-D>HdF(AV?EFZDWT<)IXG&0SEfZC@\UXf@)V^AJ(]?-/LJ\=
8XJADa99\Vc1fW2];G4Ea=a)R-2#:&1>=>@cPa8N<Y>K?A5VN->1QQD-:^VHa7O&
&=V&VL@&R[_UK8Y]@&^+O-HJe:&E6fO:>ID^J&Q)Xb:9HX^YYF1/&&4Ab)SK=902
OKBR.[a4g=Y0P:9fHKdN1]G>6P@,ZH+WRKLP]7\\T-T05\08a92O)00?;2<@&IT3
[fQIFbF6a9K7O7209()87P7L_3U^_YD3WA3M?NE]W6\)d59.3#T5d/#2aAHT_Y^L
f7]cR&)fgZ6@61>BP#TDIZ#=Xf6/b,&MCD:KB?<HCO+][cM1(#cCSb[1-GCZNJIe
RD]2JXdMa+\=7YgD/1RcW;#9+4L))L;^S.9dWgBKBK\W3+d,1QdVBL(J7E:MNWO1
83dF&NaX5ED0gH;^8e\OddT^GYgD/N?,1]TH.<4G##N<2C7B,>VDJ>a8(H)K)LM.
;<KK:_IS?34O\E4F&&;CdQ(\+N,ZR8TYX1Z0eeY@f1K681LbBR@g].>0ZYJT[bSc
H,Y:OcT?P5VLZ;YUX=HW]DcQ-,OTQS+U-X^b>D-Z>8CZVe/QG3_d(AE\[\56G4RN
(eT,R\]F7MZ+RB0JHe[SZXFG];<,9\_G2)Q,^,S&H:(S_NYBc9NT2IgNLeI)3P-]
&3c)C&]-,gZgc^]Xf?AB&#F/W_U-@b[0X#M-,9fdYaJM^^bL,b<0)a@>I58P;]cL
]]9-H#5-f9I&9GKd8/+2e,V0BMY58@B<OW/K9VH\(^LL^MN8+[S1fVF-O/S\2;<N
=M3QU_REY:JCZ)e)+JQg.(@T>><(\Rba-6)41eFHPdU6^=1Oa@A33H6YH(\.<G)O
C1]4)[ZR_Ef)_;P2:>QZ@JQ_FH+I]TA_7/3bK?-JO2\cKHU5YGH.a&0d3bf9a#W7
S3c,ebPGGVQIZDNX]94dP33a1SfQMKV\0IaX4T-6.aKdc#Be-Hf2+3e[3VKW(8VS
M?YD7NY7H-bRKMU7GV/G2S2<5IO)(>,\AO,X?H/:<e_SCN/II:_TNF]6ZVXXcgBA
Y=&;EBE)X8..PRVIV;9WQ_Z[b<J_:<=YGLFR-\VCKX@f2N:1KUFRESAS09NI>7B#
9;CH3P,6]XHFT--cOTL;g/@aK=E^cZ(gBZX=(K\cVe\-E4OFe5]<Tf9ZSM+Ef;LE
35fF=SbcdZZ-L0LcQY:0UXL:R[UMaB6P]KSYA?G=+=b\P_GGV<@:VM;WGV;0a9+:
S7R9-e)(B=)FYg>MJa6?TXQ\.gJZU5A2.3WLXb?&Q3eP(^?+N;/YP,OS9QA0-Ke3
RgKaSF>\NTO+W_ZIUZGL+(@4@Q\f,18/;S\+8f3]H][^\_[Q<3f<1=Oe1#HgU;bD
J8.DK:U(Ae<Wg?Xe5IF[NDDQQ9F)ONUdODGU5e3;IZA0&1TXO2OOHbZ+D,2>d)Ec
ZWF^#]H2]P836N:^,#ICKJG[QA;DGQJ(:84+_(5_2J(22@GdV7@Z?PO/Q2#b?AOR
EOZ3CZ[AL9F_WC\C0A69IR:7Pc+M?&0Je/G?K2RSaAKBQ&/CYDOeNIGB3.>1+JIL
VKA+]KR5\(/_T=-L\QRQW[)]#+],R3;Q7LLFCTQ\a]DW1^_dF3.Y-L:/CTBC9[+\
P[_d^01ZV,9bC#BU:G97EE1S]HULbG]28+\S\MQ?W+PVH=See=__;_d]_c?-ZXIS
R/9.#QPU80(4^9daYIJ@dO,2RdI0C<NfLQKKF56,&20>92+9(\d>af8P93TU#ZH\
QcA/ef@S7ZJeM\0](8fKT:F;Z@7LM6L&N3312Z+5X(.EAYFN66f:2UTI3CH38><9
2(CM0?#5()0c9O>0_V5;/PNSeU:G4eY+b&DV[RLgb5B+1FT5KXMa-=Z:J6f(IS3^
2f;V)09FOX-DO]d.LBK:<c=3;:IQW\D^a-0^Oc43cgEb<-.S/9]c4QI]\;8B&9Na
;=P+NB^)4UST\.T:1Tc4YP,fKU@YZ/,+bc\:MDF-0^P#.]cDU,aK<2V7cUgJ;TUc
1N#0L=WagQU(4/6[a2)ZE_PTCIROdI5_Ffd61_SID?]S^DS;VB.4Y[Z4dKE\S2cW
8-D0P<[7RN@@a\/-=D0;_bV&2(SF/C)N8<5JP\MOH=#FSU998b9:W5@;/<,DGLY1
)#^+?GLW\:XgUV\0SGGH:Cd(MVFKU@__UB\fT-bU.JO^E[b_5.Vd,5ea>ZB+WAZa
)36:Mb[9KC]J]=>50^UP&(:Y7T+/Z-4A=X]g.U7>2cNK=/0LQSYOFBWF+M2Wf<]?
N_O^8D50O^:2=PQR/-fI<SJPHP/d5O)g;R-:VJ\.W^UH^K82W:1(K4UO.dK@SC;1
96O#\1]J[H85TYX>&_M9+KNdf_fKE2Q?SQbaNC<e_141IgCW;_aR6/6#-YAeZ64M
_+]S_-RQ5S3Z_VLXNSOg<U[WXdWYb9@fYERL<4C0UR7#.J))U?8YV]acQ[BG=+F7
)#P_;#bI4).+fQ-EL8g[;Y:0Z(1dEL67OK-O]IAQf@&IGC091L-:gG7(Z11I]81:
fEJ1^YT766H:E>Z^^XT:2&91@69@8#/0N><=Pd8OLV0?CT00b17I68E&QF\&,XU^
3&&e=aQ3^X)2Q#HD8e63)ED]]M_=#@/.ga)TN?=\d^XQ.8H;H3N3_B_>e?5KHaEb
K:G85M8d]cRR8IdUb.1,(Q&D]PWC>[/;<Fd4RMRXX-D(#,.cO_AbP+ef>Td]NUIF
82g3J+PR-XaICP69fHOR+bPg#BNI3;?6@=Yd_e+2[-U\XL+-,eAW]S7D\J)>V-QA
):8_SY+V(]Df58O,fLg5JR2/G&_,DM7I<&CB@Z)#bA;?ZP.:,=5eI&QZNY4?[8V0
>RQb#\(3>PFC\B/L8.(J9&U)6fPKd8eQ?b7UE#/GV@7CX\DeZL/1D<.9TGM2-Fb1
4:?#TNK25(8T^Q8[=ZUIZKO(1S.g/C2^WL#[KAS;HI[H<[J?8.>LDX;-@BP99TM_
?HaOD:9UU3I?<.V33f@AZ)JEK);FM&<E&AcDg83+#DJ8C][c[;2@a<0_+aHQC,5@
2G[8QW_-E[?dJf&V-OBYNZM/00B#GH8&;c&C4L(:<.D-S\e9f,e;J)7g-=TcI02&
=:?cP:B8ZO4)Q@/-IeV2-?#T9R6c>I>G/5fT4>I5W^;Lf/^=;+O1.S[QfW-I5MR3
)dO:Gd/4-^M3S\NNGfUP[c=O(\[;@5TC_V_0eVYVc\44);)LROMWB3_13;3=O==L
(cNT8/L#B44LEZPV(bcIV</6X752EG(T4U<0b5H[)#bZGI2fL7AXRI]H\,+LE-??
VLBHWQ82]eWDD-3U^f3Ma8g(&VGF-Icec>2B6+9?Jd:PS37F<,QVS?^.I?=U1(LZ
VEQI+\gcZb&\?2,;AZM4=X.2DL8N8T:Z<&\g3C(CAM8dW<5T^JD?Zd+.?&F;;UEU
0gZ\IONRg^X5R\;]f\NOfFdC.\7?IM(3dV60O7Kc5DOY#JWD>9AHMGMESgXHe/]+
9,?;^gd>ZA]0N8_([WD#05(E=N3LdDBFUcQ^RH[WN?O_Wa>-UO7E?(/55GFQS,2?
DMI_b>QS)]bU2Ha/-9UFY;H,=47HP73RQRbP=ST(5Sb&0XfP8]>+F?1PIQC7J48Q
T;&E?g@5E9H7TG?,NGAYBV05_WI^1\,6aH[AM&/T=_FK-9B_=FOI/NKg]IOA3G:U
d9R-Vd6ZLI6)c<UQ^;)g(Q\-b\:>Z7W3Jg)OXSU_6PIBJT(d#&:+ILUdNOLOHUA8
4&+YU-+4&YPTAU,GX<;d5=E=9,P/E>6MW)<K^,:WPgcFFXMU:(c#N(X5;)c.FBKO
,QU\2:+=Sb=X:<Z](,>Bd=-S&W0Z&UNQ^M_e+N(O)K9-KIf>6^-I9ADN,Ibf3LXD
XM7_P6KfA.SA8HK9Y6^;/=\7cS]UDQ0+;=aDITHR.K,@KDgZ\6@L.R]MaO)V/UAW
,6099]<H;UA[9Y3#14X>,S&B(UC6Q]e-WWFWEf+UX_&:eOU317RG>.EdXRcbJ<1K
)D5R@AAGeGT,#,-2HRG@NQaARD.\VT5B\b2[_FE7cJN/IOX+F#[&0bCPH6)+Q\;C
>D]1TD0I(.UZ-f-(^B7IfB,9.bG^8R]f(a/52VTZ/^Y.A)Q^S[McW[4Tc\OL]^,3
U\V2D=g<dLQN4XVXTcXO)[NE=bXAQS\IFH2&A389X1\I^f<(1BS[&c.X,W]^EJcS
G:e9I-&Y:5HW@HY2Lf2AT_GG.H:bPAPSecRP=bQJE?_;Jf6=aR>F/aYMS>c)a4Q0
:@IPK.G[0\;3H/_M=\\)1?-I,MCZ&<=2SbW+AZF#E/aD[J>YS&<f(LE=V64];U&Z
JVN>EVJSeFg0B&d_:X\;-_R;=gc#N)4FCFQHHbZ(]e?WV_<3GT3PF+?&a0(\A#^)
8_^WD0^g5D^@RO4]-,PUS-/bbD:GI+R_R7CNT#G)IbdW#L0)J/7Gd@WQZE8A8=LI
K8YI2]O<ID;be#5^)TTEbS3\C2cI.,f<\+0_02d6Cf1X[N?H@1.D[bB0dU/Y<#&c
NR.X[&ASa]-Oe(#aTe#[@OC=^Wf;TTKc2Fc(JWDICU:49CE59fD^-e(Q4d>DCW)=
9Y?Z?J-QTI]+S8TU/@@?@MbK9QI]f?3^C2/5L5\8]/.#O&e?Yg7-BJ:3[,XJ([^1
gI_,0XaB059P&I_5C6#,40W/DMONYYeHX.5I6Q7-XKTF:3a&gf+c:B.C8T/WKNC8
?.B8]9Q@K]74@)^^DBLe>b\HVc6\cV?67cBWV+)8-0MSeC\?eAdL+CG2^>]L0S+,
82L11A#MQUb+fa/.e;+EA8,TR[I\-\?(GLdDTba5&G?0I:W8-Q./Y7<T[LQ:F]7&
_8gQQ(,Jd<:[M1J5Y6P-(Agb1FR>47Q=X>GfM#5&Qad\^a[_3@7:+[A,1T&Tgcaf
<gN0d4?K@3D7+VRge-WfJ0JUI9)6Sf)(P=12#<Z=?3E5TW+U0IXFX](4U#UE@2,G
be5gW5K2T2H?-:/A4CG^EMdA[&WB.7NSZ&UZ.;5bKKH#YINSA/47,)Z:aL]2ZagX
[de]<U_6)gN#K7U@BIBRLYF7ZH\\b_J9JO,3K0V8GNd\>1@F.Y4BbS(S7a.3gV[D
NCXOXNR\@J065<W_8fIgHT\fCDNgG4M1<#AJb]HIbQK8HG0fLGb6#gST5MdQg(Z9
OEB(;+K(YH961J2QbGJT(&YfMg28O?YO-gcNe3V[7aD02_@LX,J.&>:)X>cHbUe/
>1L?K]LTbX&&=P99##(@6/;-dL/F@50&,BcRO5/1UV.@0\5H_@,VKc=R92CO1_VO
TM-a.3I?bT-IRT0XSbP(8LHKV:Da8U=MWC0b=6A]c6LHU61-cQ0BA3Wg2F,VVAf#
D@C6@[4L+Y.YPTM1X;3G:H@0gV)Fa[O;aPd<UEbcXU@XC?9gd2<@<.fE2W?^L\g.
[P&.&HG1[JQE+/96T1=[CL[R4QO6?TASGC20ceTK49e;5LQ3W<KXT.TGG[QXaGIB
/./bbba_JH>ggdf3FGdM[W7>W2b._]20D4]86+@/787[BQ?LV>8XH/>GO;(V-FXZ
Ab8G7a:3T^+1\5dcbBA#0YY;=<9\/IX@b5C^SQGVZdG,J]F:EEbe176a<OW^;G:@
QYOUP[<eHMFHF6-SZX>f@P0RX>K^26?c#NA5C>Mc(;gZTLD4E)4[^Ne#<\ALR7Q:
OVYYGAZ.fDD>R&g\O>eS#Ma\=(M3b4T91cYEfHY>T,>fa&N39=1Q;4Y42,<-S-c6
aH896J9@c/g04II<<2SUQPK/I];TJ\NE[SL?(>;4\]Id-)3V0#/_Dc+])\c1G3:I
dP@9_9S=M4@XT/>d&[VM\GL=7)FT@D]=KIJFK?CD_&H>J/&L#&@RHbR?g27FTA?_
B&()-.7]7_OL\(+:bG=C>F4Z0N:8NN)HLX^Ca6eGN@\S1F+O@]fY+8K7dGKF\:LA
YXc.AA<E=JO46YdCYFZdXbD\4B@@C@K),0,O.]L??_2>D&;G-f#2O^DL^?Sb,:BG
OQ-P:M5EbPL9RbdJM>=\2.=IH:Q.6cIPID-g)ST+IAE7Y1DOf(KX)0A2QFd)F>LS
6H,.RG4/=f@:X+]<9S:P:H9F8fU?D[52D@gQ?+>R6=8+6>Nd#(A8J4TA/;-)=LJX
BF\;4&aQO7;IHS-O9K7I0H)TQV=eQMHX>3/5>AcD(]8LS)QM@1<(0_R_6FP\U@gc
g,(R,#JLC9J;.\LcREG40_AY0-L71M&U#93L@BD\SRFH:Y#=Q>3+UQW3/bDZ?ba?
(N.2F>d>00Y0Ub[Z72QfdO_L)F272#c#18)FQ)MMbY[>S3BK#FIYgT/:f;MA,]((
9<YK7A74_I>8=<I]0\S_SZCK=9)R@JV?USgUAJKUEW,D.[:)85S24_J])XMd&=9?
)6Q.[Y<;[]>9GV]76aZ;JWFWag>Xd^@B3RDDAg31-2<_Z>9KF+#(/@XJ<8UT#Pb1
Z39b\@9#BC=V2,Qd.9>=:)eN\S06]Q#TI-VOQHWg?BK4Ne_,KS2TMaZGK]EH<]NN
c/7?;b,MScgX/Ha1@DVY;Q@S89;BJbD077,GC]?NVEc27I-((0?ObLR_R.faT[a#
4g82>BWK(Ke,?4RL9f=VcE_OaTRDNDd0IZUVMa.PZI[&?F7KQSb:3Vf82I]6VaRH
JWH9P&\;\5fa>b_-XCAWUCSZfS\0>/e:5LJ(62&\(ReJN^F5\1cRf84PYPHdS<XD
g3D?.QOBUXF(?W.\LZ2<>Beb4G5\Q,dbRID[E5=#6IKVU-]2Q.6GcgVA2I>]+PSO
)]]]F[.G#1U[ZPU8RH22U5O1EWZPH.baAb6:KSceJ;K0\:9W/dKL>/F8RJ_#F+4.
Gg,GSg(.Z#D)C0a>>.CUXW7?GB>7=;+@,>NKB,4BH-fJKI,2/?-@4P2dY8O@9E^)
.GgCA\J#/XM-,QJ.VKfUR02OaW4AB?Ie@9O)/,7+>eY+,Kc_d0dg3:Y1NW-IV<5;
3f;=+@-H8W7Z.(J9g7[W^d_TO7593N4.S9Y-+_I;B@gXZgL+DbFc#\Y@)gZ#;(XZ
bEED;=E2:X;);eB\^9]]g>Se/.83,ad7.Za4VeB^P)eOcD-RG(MDf<M-3K/KIK.S
9d_Q+^3X>@AYQ0(2EE<,4Z6J7Q5a4UK??e<.#7e-\AR0XM=644VUFc-N=:=U^RR=
(@:=RP?H.96;##b\T8>V[gf?IF/?^6LXfgHK1NAH^H3cSI[QeAGS,de2KB85[cHS
<0UT6/UV5278_UXd3Se&f?&P&#g4P>e[Cb4:fe0O5U7?T&25=A65b]@V&.OVP_;R
DX/IbMNC7L@&&8c4=.G68<N36CWDEXJG^+6[^CE6KT48-<.8SH_XbMK#OHV9H+_U
^Zb-c-PUNY2FQ>5J,/bF=_NB/B30>S=Q+YgUR42YOQdfc5]>A(\\E.#>#Z3;GYSN
PJa@HZLC5H0T1/DZ-;cffXL01a)](eFL3HgTY\/f)I]abH7ZV0ZgU9-RNL>VZ[g&
O;a;d5M[&@BCWM<G6Y7Q:KZ/O8S:HF^U>Y;/62\M&f00&2=+A1&F9G\S9a#+M8I]
UD+:ggGN.)C=b0TKI4J?g6&33W=@2T&AXWG]0&460JUK=&3P^QN-><E246Pbe]BV
4f4[BH9+JN(.C-3<a&9,A=.:eI/16I.?,7[@UO2(DF+62VO>4F_TgaaV33_)\c\E
9&T-5BOQ^02gSeZN[d17L116JbF=)L+)@-B?]VYC+>,=SZPS;E?FU\Q9([@\W_7,
;2b=:&]WE)dfM?f5V8fGP^9e):K6dY?WD<](/0;f\^R4OZ7#3ME;D[E[faVbQ1M9
cN+A(F/Z-T_2X0cagb+6O0fH(#EXC39][g53bMIDc#MT91\<D,]Q?c?(X98I/DK]
<7eFc<Ua8KMJBX(C^8AHKVILL&GUP:dEO2LWAD5<G&.S)aS8WQTB[1W7,0e=ZJG8
)243N_[?J[(VRL-f#&B?B((&G6GQ50M_]#WWK#>>Z\9FI/1M5(^K8SLFc^O2:F3Z
Mf[b(/W#._-.G8bD[:e<S;Q#(OO#^BW50NW2/eN/L.B;D8)d;W];9UL-b.aH(8O\
^D\6Zd#+GKQV?FI877U=<>3:],F4bF^52JCH):aO0(fR=0ZTLFf^,\7/QJWA1]GD
>J\1D78Uf+BKQE=I0<G&/?,=UL]^_)C4aIZU7;gE8VT_F_Uce49A>acUc#]TVL6]
VB+a.PAR8\KIUR,BVD(3(T]D-;fQbf\BKe)S856K9C_PcH<9@3;VM0IgH;HO2Y>3
[]_Q/.IXE4T.[9A9Z1+J,=:F;0Fa0RTK+XHG5:C3@\C33\<+<0FW40+,F&c>>4CR
g8bIUCU.Xb8BYVVA@-M.[A/Kfa^9JYbZ@G2&a4YFQ+gZ8(V&S<b+BIRL)aK?,4Hc
gg\>8G]5cDHF5RPP@^H2+<:Q^DLU<6+E;Ef.CSQ&BN0FLSXYc[^77efV_0PeY4Rb
WL./Q5?=Ka/eF3O2,UF;RAG?-VgW@K[B<E>28cHE-aG:;H71G=Z+4/0Z<IGRIYA&
c4;4\FD7[.02O]^4@D;]RZAHDJC0#Z06]WJ-X7-9EB5P[J&:V=^e\C_?73DdGN^c
>7\4\>U3]PP=#N_dJ<1#\O(=Q/OK[1+X?#4L=K^=L46d.+S6fg2EQC037I=S22[S
YgOb-?/Gbc86KDFAH5?1GL_\+W/U9V,AB[Ce[HH[B=0I@3)bCJX2_TR1c(4A&,=N
(eZ2Ta3))/BDTR7(+([-aD3#WS1=f\,B(EVUJa2H(R@&HfXERFS=<IUPFZV3R@0(
N)eBL(:>3PYd;:H9)+H(J4;1W1X:HfK[VMg.IHX;A2/8K8JSX#;]_BJ\2(@?e4G<
,/M(SeB/6;dIG2MR#)b6HEY.e6Lc5PCW++N5PJ@@R?5OZdT2]d&^\L]/IU2=:c[)
#5J^6(-WdTYd4.[86JI4=BC5+=UO[cDdHDZQcJAGJ-=4:+12BVU=XNAgGT2)c[B(
A5U(d2TX_OTE3(&EJ3TYDLJAGU5;O@M7Z4UD/Tf<MOI;=,YXSZ?VM,)7@RXTKYPZ
WX<)O&2D^D(UgNTF\RZFT3?E0A9:HI?9_J)SL;<<[SUdd9XeBc+H-)/PM7J[BQ(3
JDWEHdW[g&THFcR:FcVQ)e]=OO[7GU09YO@(b-YT1HTE./@CZ[5-HT/SQg4X2fDN
0T;&N^.bC6O)Uf2JGg)KWQ+f&:Q?1ZFOYPgR^N[[]B973R4c5DU\DL8@N;:#c^b&
;VAN]&T3.YJPOO^<I<?F+T#JNX=feB/:>17F_:(08<5c&JI_IDE@^3T<8;Q-4L0M
H@.SD/)P_M8WfULAC(.XOZZ4E@W5T(CK^3g&=6-aDE8.KY<D).S@@I-5,7AHC56.
A0,AW5=W&_IT]:4:[g_):fBRLccYY.QNRB\-gP<1+&d^8VJ8,;4VZd\RNF+Y>G8C
PN9&SL@58/6X87P<Za_Jd3eg1225/;GCd<5&WQZ]ETYX\dNe)e5-.#OBQTY0)DX8
(H+D#20L[QB[3I[WfT#6IX@OP?+,XcB,P4@DRF/]MBIL.U,N(#4AL21;a]U[1&=&
,,cDEYXcdg,+H?5[/I3)#\_=MQTZc0/BCb17:0@P,2,WL;7H\dC6J4@_)J<)bZcP
5O\7KV5->^c^U(75dY2+a9_c>.:AK(d))9.1(W820ECeO+cL^O9ICa-D(fH#/1AN
Q==I\=-a^:Da08#15G(ce]__=(<C,36ONVM?A]KJ..]:aHTI(XH^@.8IgF?B(fY&
fGDZZ@D@DR<=;f5US?8?c.=:\<cG/JfNg4EBKB3MV]NVd+>]T5GZQK9DJ0cY-783
#Q4D&PKb&TU32fF#aF&1eG?MJ,OgK;ceN#?+-+\FDN:SO^AA4@>5g@Q1AF8>]U;(
Sf(^@5-6Pc\JD@g3e>4V6T,7gLSW?9fdFQ[M.&#7D8f=cfS>Y7fQGg@1MbBR8INX
XIYd4[L=Y?eO3Y>;RMc@R-&4LZ<P1Y9f2V3d7?<_?>Q1HSb,7\OYd-W\-/g:Z1N>
PDQZU^K2>2E^#JFN>a3.VCB(c3&H-\)7eVPY+L+aL]f+XY^N.Q0gH,PF9FJ6[Igc
I1d2:aS\OP7F91_CQHJ=E#,XVBf99NF;3WW<dJN=,DI)a:CQ@N<c0ZHZg]DVPcV8
KSA:RbF?H/U8U)Z8R\2=4[CB5e?M@\3;+.H;L=Fd0e/7KIY^N8eg)1[&e3)bPUTF
[0.6#LQX7a9H,>LQ>[L#-c+NNCY8)&Ge)[+e,\JU5)C:B-PdOMYaD]AMYLBQ72b4
0W5^e@E<U;-RE&4H(+LNW?9b,&L2[;&e7/F5CM,9-TPJ-EFK[d_6IC96Ybd8QG.3
c.F>LL[Hd+2b9F82>BTM^==1C)95.d>#LCKaJ57HX<T[3[P]_EO5RB#JMWGLA]2V
gG2&M#>W/8d1,PGaLJ4E&OR6_WXSeT(FNSc3Lg]CY2OJK6D.[IRR-+R3:^(]a#fg
Y##7]D7PDe0cXH#=[O(:6[XGQ/AQ)D-(bNJXH<\^6PUg/@=5HDZU1F(S,F&BV<?(
IK:4OS4OO?(<(B?(OUGIU,0EBb_K@-)eFKLNQb)DE<SVRG;TME>T8dXVF-BSAPPb
;A=:T>WJFU.\:G3bX),(/NBQIP\/4>WR^V/6=71dB1/Y)+PIaNQ;;^BO#<#X&WX#
(,7;+]?<=6?U(,+]2eWeGJ2\/DLU&:44:d<><JDNfce7aRE_\8]<>?1TBO8W:K;)
fA(SDe(6]bd_.;I]#))0U8D?cS(:IJA&=b?[9<<ZG(fRfZWd3N4+]&IBZ[,F]/d:
3>W_DPd--MLOfb0566V;&P=OEc/8R;?d#g7II?,-GZ9QAab6aYNPP5R?^^R+,2:;
N<D95g:2UO[1N)FWg6O4A7SSXg#Q6DXBN]^,XbT@B)EVf\BLcLaYZa4J6SCa7P>Q
#Q#-X6XdDXNVZ+cd#S4>-VeQW4#Z<cLDUcfBg5g_IHFJX(QF==<6N.DS@/IK69XN
(+>BOA;[Xg3\R:BB3eD(]OV.,FTe>@ccHbgZT?JJd_?,4:a8J.146#O6E?d;_(dM
f#NO\>)1FPA/b=^(7g2TUOM7R0:=R4E3I]MHIe<gbXHRc7YXS7O)_(QG,-3fTOTG
8[2W?ac6a&OJUSV,I/)@S6MQZR,_]SYN2]4OBZ&8(#dX5CXI<N;dMTO+-O2)EU?E
2-_9LX,@d8+b:14gf:;3DH@2d>)Uf2]W\MEB3437D&R.F368)aOLe9@9+Dg,VUP;
5:bDXQ4U<L--L<LgS8V)KgNA8U\^6e?cLJ=c?]6X:DcfgJWIe;aV8B3\I]-.E>C?
J,MdASFWP#W-89g:ebJAfF?0Sf)]gc[JJ(=IQZgFce@T)JI0gFWBg#Y+^6X_4J-A
H@IV&,Y&86^N_.-TG=7IH.F(b7/:@]]I>2FG?CJZ&QO_NaC)(,KJ@-<J93:]67,S
(_L:MeddWDBHBTB)J@cZR>&Q3K+:(#.(HOI8HcHZg-EX)PcQC=&eBNLQ,eT)6A55
\gWB5)Ff/cefB:a:FNU)RRY_F0_=/.;cDd]b(D.MBNBXdH3]L@JSe1H(OJBGD23J
#N7f\+GNY#(QTONF.Of)=1a=ULY^RQ7&c#^)<HP:YQAQ]+g?XOT<LgN2QU,5PHG,
:gTZ&]Z,06NBb3fC,7(b)\@Da\60fOPgQZ]@U2+#K;&)&b@19,[F1GCFSE9c3&:A
#9@>4CQC@c^f_)TPJUALXB-#&>f2QVL9Z(b;?NLa25TeE6]L&ZCHac^-R@0]TQ_V
W&0Z]^O9NB(3X:T9eV[P(VJ)5O.&X<]R?16&LAQ;IcgZYZ5I_9]WG6Bg@fB8XH81
LM=?#e)Q6Y/3J5/(C&8U(S\@OHX6^gSB;H-L<53H4Z)Y8OMNW87A&DR<a/B;bS([
dJc:2Qd37,#)>X3;O8Z^DE.R;UN&:.ZS(-,8U4VO7,=@,Q9JM>1[3gcfKdUW@HOU
2STb0H#;X5eH9VD\?0V6O#\F2T?2XXZ]XBP07.U:9G,5Zc)6-aIOO[>L@I(H4../
b?&>W:8PA4fVLa&ef_Kg6H]XTeCG#8e.,dC\\A\JC\aUKJYFJ,L65(K218-7K6D/
Ec@_NM&feAI/+/[NO->6P?&<8@.@dPUQBFQ7<#f2UNQCB4dYS.bX?^2g=Q/?N&+8
^RU#QA(G;6)GBH.(P9<&XJ)Hf)b),f?)&94G_2]CC@?+@,WE,YV;aN8\;PA7O;G,
)Z]NFVaZ?L8BgXUQ9;C=NMPK1=GOJKI2Sb8_Ic3)gZC\1+ULg][d?=&Tc>&c#H9Y
8ATX.APcX[c+T?JTIG;_Z+I1fK.c[XfOWP>@b]@9/(Y?^^;XP4fEDT@=>g::f#+F
VFa<S3X9V6d:fg/O,3XB;FR?872\:0#ReOg4HdDXUBZNPQ+J(BUfd\be7W@e-TdX
-,+2D0Y:E4WV]Oag4U(/8D-D1LC1fd6MMVKXa\;H16RXNF=^d_=V\?UYM#03)X)8
PJ<dGA:ed>@=1fRKSM7I9P\e1DV]+R_:0XWFM1:+<R<c[X&1P[a)W,Q)62/M/JVY
[ZB5]e(GH>1PIX\/8YM43NTIV8+J0eb9X5B(/2J0eF&11L,:-<^(FB___\CD-3N@
c#W7Z^7<,C>g[_:]0T0W27)89A<.Bd9/HH9e0O;eE;D733+V7+;eGNE-g]VX>MQ3
B1LF\YMEV88J<3KWSY<T8:5/&3S.fV9C&#=(?g:QCS?6@SCBEZR+)Q=,N&_gMbUK
eGaVZa5O)ES=8;82_NOb<[HM8\(@g9)5Y&N5N/O_O=F+eF?K>UB+8D^QSaOTS</7
M.7J<=:@J4/)8O0b1BDR:BP[BG1?H#MM;f,6c)4KJKGD/:G1)]]E;,C<b\IJIJQ8
c+GUPg(f0MYV(-D_f]AbK(cXLX@Z:[,<M]I8,eG;4)Y#PbJ#7Q48<Dd)R\&9,D4-
g/FV#2Od&d8;EO_WE.4Z.E5GCQ/BUR;#LX?_ML3ZVUd?Yf3?77=1A;.K7ZGLc^?P
=PDcM+Ic]RB=VA^H^IF\MKETBO:d>/_HWLYI1eK&aEN:ZLZ@XXX[X:#W34P4]P3:
+_QF:ZOaP(67d_G+J@c-\M.8#Z4L4Te6<a4K:fF@Sc26b+_eG[9QVHEKQ)GNIg/-
8.6e]K.6_F8#UDTM1-(=<:]S(eG<ZX<15^XegCP9W+eB..]YbPN?af25L,?SSQT#
@0#c9WIRed=#/g;HVP]V6f+;AW#K41R_?IfTc06EQGLV>EY1+H;.E/=.Q^/ZP_OZ
&ZP@>ba[VTC,I(7[?M(-PV/#J18fcG25+C:0TC=D#J,,AHfb2)Id&/Md@(TOP97@
CCa^-JX#XQ7WfQ6QcfX/9.bcBL4_G>2I?8,0G2NC4US\eGG\Y8.=HgB>4MO)8LM\
O9Z3SE&]92;[-gC&N07aRF?M?eeO4Fa5Qf0cXXa[_H8+EXLHbWO911W)C@33G.,,
3>JKg7:=bb#O]S^?GO04-+G0I5Q3?=COD<^fW;3-YXXIc5#]:XfKQeIZ[)]gN6C9
J:E61E0.Gb?H?TNXTZBI9FP?\R3[0J;P/]()\=G^0D5_P8gX0FC\8(^M\d^FP1,>
a\AGF;=G/^HZ=P5?CbT:VG7EYLN2U_B#6;6QR-U50+).P)=9d#RaW6]/gLX=Z=BJ
&g50GcUV\WB.[M.[J\LT0[WXSD&GE5E72WV_=XF(9M1=A<?BB1PPGZMXdK(Ra]UV
J/MG\N6caQeSBdf9bC@R77=7SLf&I;,>GRb)D2[,a((F#6\4_3E0V)31K,5N\8.#
NddD8GK-S+R=B:YAE(I-SadW6JH,XYQ1<H.fIPAS^?Ag:)\e((\<E.PMOe?:PT;0
dLEC9-VU#>K)E3d\;b(3?0O@+?[:(2._)-IW4<V2,[\&RW8G]K3U.0(60[f4RGI2
<JD>2#f7fR9JI8_>_8OSgX+\PfB,6g4=KF(+Y98JWT&UUa24-37FcL<T6OX3ME&A
AS><+IPAM6-GVW]+HRQFL1A9S0,X-0P<VB7M,8R@AJS<ebVSO8[[-1?5CJ;>/TC0
BJ7#VH\,A#c9B=3#S15]DWZU)TJ)T&F\)]&9?NSdUZZL4KgCY.RL7EIO)6BN_&];
;(Y4\WdM=.UX[#;N@LgUQ>S&UU0M^1W\5GVbO+?@D.H]GdK23\O^]7e/:@:].P(N
Yf-.QdTQS[XT;4)-g.T;,R_7W^I>SK<^Dg3@7=.2M8D@]fGdMR\6#0]c@2b+6AG(
\GOO#Pe;4[b^,@W5c5fWZZ^L7^)39QROfHU-fd/?eYVPe2)83=K,.MQ]2I1cCT+3
TV-D<YP_5:<,9TKZ0?G)P,IP1M]6\6A)<?Z^Q,<//LKf@]MDEI;&gbYc3/GTBLZg
-a,8e<NH8<_-e4[]WD\gf;AE1C<df_6)-7&_Z^F32>C4Kc9&8AND_]Z2<Y<AfC6F
;I@/0TQ)^H\-V;CCe(^6Je7W9QDbdeZ\^YT5Z[]&60)&_=VCM9Zg[(C[2A19bV8.
#&D1f(.eg.TU#E8M@^+CEONdZEM_S6IL^:Q(a@2//B8bX=.5VKY_YKK0[,/e+IDX
NS33V0)?F5g+eII[A(HOd&O5f0VBDRP?D10^@a@9V_f>N0NLH\3M2K:W_K;FbO)@
@S;H64d[/C(C^=RXBUTM-TO6#::;BL17ddUCBQ[X)0F,?IQc4XBH[LY7f:[Zg8M7
g]EMTF\RE(M_HCNRDPf[A^7d4cZE#TG#^MW._9MG?38)-QN]:\3J^g(>PS;D4M>W
KNGJaZ8@^1791&eFL>A5&HFTTX5O1YS7)Cd(2ff(>U2EW-3PTIT7a),8BR(+3Be#
^7<[R8UM)+4&>7R>b]CKFb,bcbc)]WU[1VK?\A=N)GX4NS2UKWgITcHTQe-XGD5&
0K0@Xc;VR04YL5LgK6JNAT,LOUSGK<2TbDQ]:FF.,Z(&2Kf]]F-LY[J2:J7L4IA(
KC;b7?eT5.D7C1[Gaf20;S?V\U,A,\O96JG6Ea-#9E=@^A6;H2?I#5:KEBB494UU
;D=(f^(5O9-:O7[Febb)Q(AAWID,G@NJN]_<K3EB3FeT2ggN10;5Yf,=J4BUPd8B
;@R_6>N4-B>[5R_3PL.+9#c_BBe<8I6OR=a9FbNMgU1f>BM.5DU7(+A\_GH10aL_
#d&(OSg=YEO9b#33aFL)U4\=#M01VeJR1LYAU.&O4c\UDG#IbM-7?4Y6-d-K8EYF
c-UWQ4+3U;Y=L(4^egF(T=a[1a;3NXSS[RA=d9a?1<.Y_/)DZZ)=ZU3242W55/C0
20dCg+&KX6_,Z,Y:6gf^ARIHUXFJ-&MV;.RJ^23;\3b:L:9V&)YYY,HZ5VKTQLbd
H3[IW)&[^4.MH-(@YdWSF<5AgG_EXBWI55@)L(c]U)YgTH2fYc18XEEDW5EdYK_d
F_eJY_2O\eeL\a.O)d0Y6cR5QNJd(b)b;OAV.5.-8F3<R3OXG3)ZKNFUXCHc?/F-
CW5BYX^3QW@4,\a?K]1c(@S-0dc+NI&U/WV-b++5[4(F)&MG_=PK;VCG7O55IEX>
/cH]6,OefdZA&8JG=Wg31;)OA]FZ.6W+H,b0ZD0FIYcRPUA7@3FVLgRa-2LB/Kc.
I.-Ic];7SSC9?gURaL.5)9RFNR>fZYfaDfX=PPN:/DNUf(<)-4KB@K8R5?JSF,HR
FG2,R3#S^K>>EYZ)YWPP8dOIB853eLLC4:C6+3_f[BEMe@P,C_C\3eaISU04(3d+
\3N?FJJMN<DfUEHLFNG^KBfJV.N>V5-AMS94g)Zb2gS)e1@J@[RYR:7AR-)<MZXI
7+ce=fcU#U#^MBHdZH]\8DEfYI23=[S,QM.R,/H,Of]?IG@:H5F-KVe)e;KJ7KfE
WAB-GW6g?J+aB3DR/OUgO.Dde8e#0Te]?W/W[4@AS\NH^H5?6^K#B-J6FIYD0&J6
J.JUd]E0+])A_>H^HaK1T7G2:Sa_\9/M#8/=]ARgBE?ITCb]HR5I3X:[V;9LG3JF
@E8CeL>5)GEB(1F#b1C,P].8#D<+11DW+-eD/I]Cf;];6O_7bPTU3QfMYa+NIa2A
\_Y4=,@&-+U1.B<X&JLEO+UaV?.;=0LA,2ee\Y^LbIgfL8H6VSZ.P;&edZFUS_00
La6gSF+:WE9&FKMBAL]\f2G1KJB&V;+eTK;#^c):.?7ZUDZS6fg.7PQg)H>WZbRV
a@e[8W@N-C3B)V=VB.#P05aeGHK>^9VBbXQ7=<]cVA\.0c#?>B4[.UYL\E8+0)ZE
4JLESCOV,5+eORD8Y),>f\\1&#FeA0]7Xe5W2INUf^RHX3+&L[6>PR@\R.d<>NU@
a/=g3V&8S7e?BYXY1&HJGW2L@8GZOZ=1))_>N;T+DLKA2S#_X9UH)VV53;^9>6(f
WfOQbKH7fT5PEF8)G+V(;7HR<W&_YAJZ]4UYS-fQfM;:XK\T.D1^Ae7P^8K<RObS
R30-X.][5BXS:MTCdQ7+F6bb97-Fc[\g+X<e(+O_2MIED><>:TLDSX-6(^6IN(/c
HNd6X^3PbC-Bd2C#,9<U31]GcY02:^7d=NJ^HAa<^R9<dFHZM97[ZH)MM<B?4>aJ
a^;5Y31c=L:(/6GRRE6CB)a<HbCe;aN,_ecdT+?gYg9(2XSR3QAI9QYbcT(A?R_H
PI@bR.MG7QMBE,IIS],\GF[+D9P8+A[H2.[OK[E&85@GEB/K5Bc9AQOFK&(7:T^b
ZX#X79),Q4>7\7aHUC?PbXbO>F&\UCN&[W)G-Q[)(H6(@?/K6E0BB74GcCK@U&EV
7<.c>NT5_XcGE@^GN)^NZbg342Wg0&F&.U1XQP+3.T;PTTOV9.?-^1Z]H?\aSa9@
@>KSXC_gJPDB/a+=4MGg]H]-3edX[L5+(5NUP<,<G:S(FT<(dMC0E8+@Q0#V4W/E
EKd[9&(#760L5]e-V0PdgKNW-1&O&YNb8IH>[ZDFe81(KT.C4+^@:^aC:(3cT\/N
.\B_76FUJE&fMYN,OH\bB_4^[eCB2G&8?B\WR77AL(](RAZc@(a<(aA?WDFI6aaA
W(TJS.>+O]ABLC\9=@6#NJU],2b\LR[,M-Y\FBU/8=E;dZ.N@gT5&J)E#Z5c</d>
.ARa#ddGFA/,=,G:@P0NK-+N^M=g?>:>IQ9/U>5Z4HP5a;,gHAaIXI?>?,c[^DJ6
/#f-@:]XH)H?8dQ6.1HMJ))3[VB@F>8B)7X@fZ?<3]/JXaEE@]GgV<3EVN5:3:Ec
OZPePXZ=D-[K#gIFO<NWVg4XAb4WNR5NM.QKZc<33N)AKJCK;0W<&QTMR#Md/TCd
?^Kf^51?=2GZF3KBeTLV,0P/HMF2\&:_A<1Zg_KYZ93)TGG)X/&#O)7=7Ra\EHO+
E5&SX1@L&9\\>I>Z)BA@.CN:B])NG3gN+W36F1Q,_gT9@Gd.WC;+]f;VP+ICJdaH
=P5F\31e^eDaCN1C4e7GFTT_25=.9(9B,QGZd;80C_0C97_1#fM1f-^WP)F>K=fL
R:_NLa>8fJ8T7cE,CRX?OCJ5C+C&STYMd1[H\R8KgUBZ)\,3&&-H>X)g;>,M17;9
#ZCG.E#W7a@XL<.?G^LgI^LY[E=?5U=MA(F9?RP=/:5eg9I:4RRc@Fe9^W<8P>&/
OJfG#HIbVM=W<]81Z_RL<J,;/B8M?,,JeZ-2A3D)>VH4=-GCR[MSB0BI;EGAV_++
(MAC:XMfQA2[TR&IX#fSIRN5-CcINQZE_97?7:8>.]W#Od.b1N3,=CEMg8C?JCdI
IDMBTBfHM(\Q/#0g.5gHBQJ:2O><[&7,EPJ60F>(>=X;B]^:[^6?VCd./:VSUFR0
_Q@_SI],5B\HD1bOMGe[;RPQRD-ca7MYD:)JdG5]QOIFJ<VZ;J7aaUC\88THHI(:
K(IFIDdDSG2XMRF^f,V=1(;D<BE(cO,>=_-H?e60YE=PW8f_e7\G6(DM27>SM0WF
B,#_Q;>1\GWH2<dGI-U<4HIW:M&2XgB<0F@MYIY]M(?=V>N0(AMY]G_bK(^+,K(I
2J;=.4WC-C2;Q.e4AcT.RW2.ZVFfLUZ+Y)+dO=ddb\=2/0?2daUU,2GQ9XbTUUEK
W[[b1?/X^>?GQOQ)O9E.0LKa8Re7]^WF.Ua)2O^DMb;S^.ZaR.GI4C]Lfb6W:4GF
>XJDL?LVG4;2EHH8_\JD?.CBAd]E3YZWRIMSLKN^fY_-._7?7,N5T>6A;&:\0B)b
N4_8RA1X]^L9UZH<NC=4]HLAcNT+0K2#Ce3(\D\G1DAfMd]];M,SE7KIB>eIG>N+
.I1D[.F@F-50O3]J=gF:5P1QN93>3T6#c1Fb[0\+>cX\Bc&)Hb[cO=8YcaTJ#+Sf
UWSgee@_d6O4WeU]>aKP>2]+ACCd2MX^>74=b,2Ff3^a.TRHR:XGF?_NQH0J4f?Y
->ES(CeE#T2TdN/\UfD>eT;#=c<H/0UE_(MZ].a,<f4/@E.:8^/U8DV,L/T<L+-J
)1b-GC&7::XV)[ZQf2G/]98=_FZ\HJP)XI5KG[C>c84_:fDbKEL_M(&F]4U]VL@g
E,feGCE[SM3b\7=L>OGNZ/#E4H1>-9@EE@JHV2?6c08VB@H[[AB4)??KZ06Y5MX)
Nc<?:SCSZeY_:BUF:aXSgF-JSF&Lf0Y?-6#gG>,]F4_(P^f/9ZTUf_JccT)\@BJT
,7Ea\NPJJMDH-8X2KL4]HAc;;c/L5#a+4NX-X7.7?QF]K6OUX8g5cZ9@1>.18U9+
GBeIA40SJO;R/3U4c,W@PfV@YR/fVV>W+Af?QY_4>8\LSD7WK<<bJU>T,663J\EQ
dQ^^SKW@N7.P].-X.00SeD)<e82LfX^=A(:\0/9A_F<M)MEcD5=;LeG&^Wd+f(1Z
E=g;+;.[#Xa[&9]]e<7^^<CLVe/TG_U71>5&2C?dR_:&W8gAaFD@S>B&N1a_O3Z)
fN.-2ZE,GUQIRKfWP@B3G6,8_;^e;@4+0#L8I^3QK^55cFgRD<+dH84;RQb+b4XC
f)/:W>,_KIRKQJR_-HP);[Se5?CfH</76ce0[bI]eB1E+fG&8LV4#K,K3/B8&aFH
B8-fKdTC,]Z-T_=B9)T3L+.#f\F,&.&UI&b;PEXd#U7+4e1)Q-I_?TPNf@d2X+K\
U\N1>CZAaUgKB:f-2S6Xg>5_]RQEQaK.4(fB)&cK0A(D#_4Y;TTfg34V#PBeU<F<
d-c/9P\V5YL873&=](@c3PQAAa=+TMF[Z\M.@T^PH<#DUS2LVbKN)]bJD17X?/U.
WJaa2d@)S>-S8Eb;EG:.M)O6+;O]Z,-0F^JLddS5-81OcYN-)?^:=eA/VFaW19Z=
aH9VMFGI1XGDMQOAU.7Z(J2GQIa(_;,C<J-C2Y]e[JGWTREdX1R_4GP9/Y.WFP=^
g5E6bIDDeFIT?LJb[-5@TG5UD]ZLEX(>O+#Z=Je?ZgT@E]?BaLVGB-gD8X3;P](G
58@V6)8K\Z6FaDMcT7@QNMQ4c2Z>5_b]fO<B8TU[M>@F:D&X_)K8dLD7H10Q7R97
K?;7O,KQ,;MVJ]\c&D@AU3162((6OPC\_X]cY&?OO@JF08AI7a?FL\7V21Y-H21g
#4+\(2BaZAVYW9/g-D<2G)M4Pd(@]+XDHFc(C]a2=U(LY?QTBZV@96Z6@^5H@Da=
\NA0/33ac5OcA6@>#XCg.:Q5eS<F0_g+2>N3.]PT]P]A#0bL^FO9G(Y9X;J_EM(^
@.NJ4Y^U?-J/^Tf(d=#N/0JC>9J)LBY^&_c9[3<6CM[_]@VVdQ(7P_N+R9)M>MF6
KHdILB-/H]:SVaef^f7C9VDWW?d<K(_F(,QY@#[FCMf,XRTM@E#)deQK#UL>T[N4
7c235Ba>(^P2W#@8ZY-CX6@D\cA-TLR9:1/g3ETaV^460+=]_dTEEF=&43-gM=K-
eW^4b^3/e.VHARgRO5QJeXQW5?F4]7?dg?_RH./K5\#G;U<gE2_IW0\NLO],=0XP
SCO^MW+cDB_ZHMTRbZM;X#I(43;W+VQMVL9Oc\G5-&;Va7LV=fGAXF-\JfP:SaSR
T:#AeWa99Cg8Q@399]2/A(@[+NZ0+X5E#KV,5\Wba+UXI^+C5?N6R6.2LUEJV0Z9
X(>AU4+R21&XOg4:W>Z[3dg(I;JJc=\/_>AQccGeX)MB@g2Q+D1f,5-J+),1+Z&K
1W30F)bYMNHPUO@b>5.-NE0S/+>6R/[g]Y[@<V7TZ5cbD]USb=,@/C,JB&?9A@0+
9=7-AZ\gWU2+K,37KUJ3OCN;T\]DSFcZ+cX26/]Q=gf^P2b1DSDNSCY<@dZD^@-_
eG54(Lb69V,&5DLUEO-A>QB]96HS\5agb5]TcDJBKXZBf>K:cB:7>U?-V85O#+bX
YGN(bNP<fgZ?)VIg/Dg?D55T<,Q\1PD;J_.&2+]ZZ?b0g/3a4X7_B/J;OT@&)03<
[JEVb+.0O2gO4f+0DMUG6Sa?7+\I./_9\#H4E[75#5)\8;??aSOc7T+A#GMed1D)
N\8Z+O(_3=Of7+5\&[U#>F-N6F0RUI^I&MQD8(J=<((LN46Wb?0g6gXD=2.gO4-2
<WT7+;eNSg6GU^)T^HEY55;4D)MX-##Fcdf2]W&V)Ua7YeUC+ZZP_c00GdI<-C]P
H\e>IWC=>XHGSPUE?\KDXA]JSaK)P)4S7D(?PTB+WH43_9G4ePJ</S^?[CS4\=95
Q[^IAJ?ZcF3=Y[cY:C7S(W#VcFT7CfKO))8]f9T)0EHB(/>O#@VWUJ61K2YdEe>)
J6G60c@E)c]33V(bgO31Bdd_#&IM84D9WD@3d19^4EKAaP[_\/4JBMAYc-)7g#HK
MC+P^I9,1deVBc)g6WNC6e90VEWM-T.^BLKLE>DF&X\<f#cP63BD)#E9cX@4PN/N
b-I0Z1c3gQO8M8+g,BIN^Q<aYXT7X:LZZ)Hcc5+_T8]@.H)3XA>\aVYdI]?dNC6K
Wf-.Q0#7)6^FWB7..E;3.+2[2R]Dg)Y+Z)9-#4:&6SHO^L^#9[),IC.=Wf3F#@6g
F,>LYO@PVcgGg[:0Z+K0QWYX,RK#0J:FD@RaEJL+_XQ-0;7\Wf-9M&Ree:(gOQgZ
3@:C8SbeAK2KDFRE;;.N30;,S4W<E2VE<3:]d75e3O&))WUQYHK@P;Faa4G-4]c2
6-&TeafWZT<Z)_BgK+.0\EO,/d<2XAOMY6EBW:[\J1;gY7UY,4#JZ0_?<7]QD0?Q
IYfcE68EJDRX>H^K?/^3J5>:4E^+Ce4:DgKbK/cN80fNI2#.6)G^UE^&W(W/Mc20
C=KH5g+J7A:00cY9Z,S-fU4BG^QX]TS/+PH>_40SY7I:EB+_=U1]0Za#O2(K)3UF
QKb30&>3L.UV&-EHfGTaEe4G735?=b>M7?aBR?2.:-NF9@bOeL:)11<R\?ZD4C0#
E_NC\0VMQDfH#R2C<<LSZbHM<)W3O5b[P&L2DbK?CZ](^F\TZU,Z^1LSKD@&;55M
\L&T_1J37Sg^QSA(N[;AecB=<D<a;-=8/=Tf\[#eORM4&WG#/E4@?/f6=]#ee\GL
9b>\(XQeXC7O+-<VP8(EHM?dBY]c4(E^B_)Q7-HB<XgB\UIVOGPg4UbR5?80T/3=
fDY=]3P10>T\G(68fA,,11TY>KV2S+#dXBZ\-d6:AgHX^_2d::2d\Oee9\K]^>@G
LMS6HV^(8dAG#5-2^Lf7?L(PLNKUNO4e_8#X@O>(_[<E(/;PI@CG^JKZ#5<<DOWK
I=:C_M(ACI;IS2VAU#[]bN:6\(b]CZ326K>E(e0e;b]SG1dEIIdSGZLEd]e#cU_^
MI=L8ZgQ+Y09RKCLOgG,5_a#/^[&?VJ=+@e5J6(=8KNe)0>[AR#AO[FZ@2=2]TW3
:3=dVVROe&VO0<^VcS.D^S5_Vf#)0JV\H^S[H1SbFTa/54.Y4eB@]W)_3KG<LOYL
:9gaCcdR]Y_SRD25dZd#,O\6;_WE,7-P@5HP\\;=\RQ2(K+J,1V9VTMHG(43?gd)
gE&<^]I()FS=1Z34+bZ^Y>EC\6WLf9b+8@M8BaaZd^)<:(.7+RZ^NIbZ,6]/+;1O
Y@EVA/G?.Ed(Xd&E1deT)XX>HX3]W4>2a<??<O<W-;3G[LY1#[>TX?&UVFSO5?cC
,)gZII_SC3>S3K#H@b@A^TDg=0gWV+1,\IWA_J.c/(&FF78&QN3fZd7V[BFHQ6_^
SXJ&VU>H2a=6O8U@[_E9(A&M/(/UECQD-WfB<@ef,US51Ld/VBTG33ZN\C;^.0Zb
e^Df]LBQGFC5-F(S]J4d&FP5\ZIFAb+L/[a._N];_I\IUU?&KKF7O^6Y)?[-\=g0
.3(_cC?(\?B)fDcJgdZJWH2I3]MK6LLPRFUP1>T([\/3c)N-/a.F@XdUVZWU+e(#
L([ScHU@TG>0)<f<WON#eXK@X#A)1G4U@QG+d2W\L,-C->Sb>[^f_01[95OI,ZIM
Q=+SNQ@AW+7-f&J/<dWa&O5[_cUBA;TL:@IAB2?b+/HTd^0M&X;0NN+eRD0X=0]R
)c?f#B]:^&7a7@bYdcfRc@]R0H6#L[[/XI^<Z>N^>P(@/YC&OSPMT]NPOCS?R4X&
BNe>eV?P.S+=6Ug=DOM<=;d/M1Z)S:;AEDIU/_3&c(/g8VSSeKD[#><6,2EaJ2,;
d&\=WF]H>0>UA0J;DXM+?=272AIH1>H][fBR\W-U)WR1b72K/3Y,D=#I#Se(]8/1
3CNALXNa,L-J@7W5R1EKXa?\=F\4)-R)HE4WW@G_?_G1+aD#?^^gO0V@E&)153T7
Z&@\0A3LC:ASg+bYZDVfUfBQB2eW<<A#]G]P7AN,-d?VR3S3@XbS,T_&@D,Ba(E4
Qc:fFfY)P44JWO.8)7:;g#8G9;-,:7T@7;U).S=M?@^,?,)2-7?1N2ec]U-S8TV?
^b(4;XQWf?7BV@X(CQ3>04Y_(d\7I\8=fc68@;da>3A</+N_K1Z:HOREPC[_K>-+
[@>QHYgU\#/J+Q)L^1WY@I-QQ:f[(c]\BVUTP[;a1HIR\f5AYST,aY,-F&Q7IL3P
aC@<K0TTGf9Ga=->6[X-9JGJ?[X6:aD@F(bV2@FL=:Qg?3S.S];OecJUJN8@KZ>2
.I]F8;e2?D6>4=KeQ5H^?WFW<)1(g8ff\2ST[fVYCQaa)F)\<R1_NQ]@?dbOL?]@
dPKaD2(OHb./)#)N@c+Tf6<O&W#,CKQEH1<e&&.3@C\#CP)Q[R5TNAOWMDCPG^cZ
\a6;7YAWB:OZZ2:ZYfUV#HB&C7.dY[HZ<<bY_f7;cCR6;V5gc<Q;QdSUIQJ[KQ?#
GKOE)T<N>YO\UGS<54;\85W,6BBCO.-<O,ZXc:9;ATQSG;>3gE10,b8DU_1ET0&g
H=I_9LNc/)c[bO\=YDK+^(N^U5XVG18OM1Z.+J<g1dA81GaD.QL0VT7D9&X:H4K0
8(^>dB[&((TQ.1GC^D(8AY#1ePaTZ?CM^8\-@4a@13d=#+JfXP+3[(<bWC=e-+4U
YF2S]A.Re)aQZ]NH0&OZ4G<J9I1[C3#MbVDP39S=[LYc3.\X(-):4J,<TU@a3I@R
XMIL/](\:Q+R:4C;\DD8+?/fGZ:MO+GDU+Y_X68<1<A+1V2\Y6KHXYVJIVJV[IMN
aO0_O@Q7^Jad(ZE,,11=PPg:.I__g<+^G=0JLANL(\J[C+C#>c;g[OdO<Sef0a.)
)L19c+IX#/N#YL1[@V83K0;SF/@11eJb_3[PJ3U5fQ)FZ9-)JLYg6g8K2X.FM8UA
eM1dCZRd(#^5[+Y39:V(:/bU7W4?#G+>[eM;)N_--2N=_WA<VFF>bEga>V,FfJ3B
2+IN73QP<Z/G[O[KN7ELL:F2VcX5dE72.8CL@2a@:9IWQHRAKeN9X/+@?[;G0+A.
&Kd)A,#GgKP=:9FNM+C.EBc#gVE7D<_5H?42a.IW1CX2Qcd9\F1E-40Mc6/QB[Z>
OIbT#g(RPG[TU/WJMG2c4P)Y>?;&&+9e6B@b5.d)6;FH[NOZP>@-^>//d,cT[;<H
?1>B_]a^Fg4I=&4ON5C7GIGLE,(:1?>)DMT;@L5U5c_(>G0[8#GMG6\1eLf=\3]5
ZOUg^cTfeXYe-Q<_b+\;gb1@df:Z(aBMN;b++CI639NH[-<:L.691U[c2YY;MEKL
GR,<33?Nef<WfG#-AcMHPDQ\HN/7L<d+SGF[=b&I@DK<+&&f\:T>KY<:[I/6XFO\
5CL6OEFZ^DLgH8=>G:I#g(A@:;aR8ZWDSL^?@?/FDbg#V#001>2A^NXCaL?]O23#
_95YGQ^RN]aBQ,[aH2J((U^)H/:;=?1_VV1.R-<Hf_>XPPcNCaR6)MDNa>c[+d6L
&U+eBP0YHPZ5FN)b-W6K@D/XA;[cP,/MbfJIMC1]?#_/&VMV[Ec&/Z@K-3W/+bLF
/U;#K#Ta)_9VNeUE&LPAF@Q?8NRgL_:0K5]/DS(A2&2@YWOH<cGXSMDQ;L+;QG+g
;D09Ue<>E_8ZBUY/AZ@W3VH5K8V)d\g:2cH@e7e+@)43I&,5.?XaKERL7M>Zc[QQ
4(+->213[OE&6cJcbF8/Q?18bU:HG8I/\./0GFfP9bH=^A6X[?TZ0P;TZX;-HRAO
:9Pd^TP+gBY8J<X=BSS170cW\2T(\ZA[2Kc2BWV&LO8fD9g6IE>2XfKd\&FRSGV^
#OPO3aO[P7ZC;B:S4eQ\^3D.,f:;Pc9TYQ#S)/e/J<T_ZEKbQBS9VbJd+^3c75Kd
WPS7757_d2X[PCY10QY1A]E/da(b-V(63RS[G6Y,7Lab.0/)AC^&EMR2.Xc2ZZ9b
3;dZ5+V]9;N3@SZ^aB0f;#)gZDC>8+76#3Wf<[><UOg4]U=IKQ)6=/.1I//+T.f>
H[:4DX?D-JTT>_1f&7X6M].FEaI]<WaXbM^C==&5<1;#N&FO39Ya_JaISZ>&-DA2
A[d1;_>.#7A\P->+A6RS?6^6D+3K^a9I<PBfZ;C3\3a/Q\aX\g.UEG2V#[b;Yd#R
+?2C;QMB+9(S;C&<.:9Sf(.=&V7J@5)bA[B@LdJeb=V::-XJeJ-JE<GN-D/LV9fH
=16<ILR6g1F/Ue7Ig1f71dPVBYZ?R1&BfTg_](=+.WUBS0M6(TG9cLM]CA0ERK>6
RgA0)/6TY)W=P(VFF)<Qfg^THQ8FLB.R,<bG]=CV&VK8a8+(S<,?T<+B+F;O73,M
g4KG\5NL_=E+3@fb1M?Nf7:Y:c[Id=XHD@KL#?;adU5WJ3G1+G,N&GXK)EQ)V=Gd
3@T0HcWYWc6\<Z-Fc=J[K_L_<dK_50RH9;Q3b#SIC-7aa&+._B,7EF728+]C(<(L
;W]A.9_QV5+,5XBNZ<N4@0>SeCJ@8A1O:d)b-b#]OB].F9RQ<gC22]U[)X&)-d69
W5&GQAF2)e@UVDa8[JGdeNXM-bc=))\WW;-\XaLY+/XFZd[0<99a3Cf)K_4f#W:M
91M?:D+4;99,H&7AGGS+_208#J0)]IE4&S7LOaE2MPN:&fL,U2MMgIM]E;<EE1QC
B:/F-AOWN_a.I,A3RGf/U>=XCf49F<3XT1CR]aZ?56/f_Nf/-cO,846TcL\gdN._
L[J(KPBSNfK<BI5;^,/>.YGJ#\&-_&1GZ2EQc-PDSX?CA:0N61OQ;RQ=F6a<F2IT
d\45P9+N.RP/aRIFW@^?@FK=9D+IgcE/SeD:&4TUgaZ2GM_d>RNKJY:9+^3=U-2#
Y3>bAV\#OZdM;F?\#+NW.RN-<+8(V&@G1L:Z2,UT)37aVM]0Ge-1CDG99#,a:&G0
c@cd\A>df^.I)+c+Y9Q/0U(8/Q_XRFEVTGXgUPX??&.;F>,B1^+&4J]TBd^8,JK,
[Qe)>:b[-(:4.=Qaf1S<Y^&K_7c:4+VA8#,.X9A?//b1Jb[eSW(LJHD(S#S<.,a@
TA4W]NK^.R0+fg[U&;#Necb#P[JPQe1_9.Z?=BK2>>[(T[XN>6/N=2Q/(KN]/U.Z
@[O.K\ZBG__J&g/aD55J4[(/.G1aS0[#9-]R\f6Y\e8cC,L[7,dV91g^UI9d5)8N
CbJJ\>cMFM&KEMGY:,R&[X:G&eG/NE3O6Sb-C\MG6L-8Q^6L/]H.LU2gSR?1/dBG
@T@-7cE]8?(I\/A[JO_))GQ0eS1IYdYQ/Y_Q<+bLX>f<BKWW-=GKEYCA[P_I\RG>
?FVCE)D3ecRG2XeBYL_6;-L/:aDZJ-96Vb_bQ\1)fLTBb1&R4QWP4V:8SEgWJ8-]
d1__#+M8AP1W4NP@FJL/QWZR9.CG^P6&)>H27E2Q_.Mf?V1\#I;.1OgUJL=&I_5D
d,O(dC74:^<))S_JdA]<:3E1VgH9UW(V98H))5^PfDT8R=(<TeT;T;IgLM/?,_6-
N;YS+)^;a.UNaQd6):c7X(c3\&M;AY\9b/8PQXaHU?a3/TY0,:E,+f=fVCL3X&JT
K+d,]cb@]d@SK/(]>9fPPFDVJ/[I25f;GbKETFB?&G7NO7?,7E;C/)7CG_3PJ+?D
-b+^P&3JeTDV#FEXcabZ1Zb6THH<#0:\+N-O[d/Uc.fM0#N\c23cPT+M_g^@QDLY
NLK1&2RZA,75ED5+A9+K5[V8F/K>dK)+Xf?>Z8,.Rg/Ng2>3]CGKY>UeGFZFXE+Y
=TYI&c5(]S?(+b4?D]0&N#3aV.A:=?a/22YLS5cNHaORU:MJ6bV9#8Q?[I/ed)]U
I11GD(a>L^a_)#EgSKD<)>GX<YRQ)fI4Xa6Y1OR@dJ6b^I1YOGKYO(3TSBL<DQ0O
aBJ+PM22,.adLa^=5I?9\)9K9?OX\2eRG6&S4[D,)Z^(.E-)J_Kf4\TN0RGcda<>
bXMf/2)^20:RD)\AP7?J\&Z><S[[EE?<[M-F;65O<aVUcfX0V(Z+g;:AH6WH[<29
Z2g=g9.d,:\eFAX#891LUZ/bB6VT^U0A-OHV+_dP3=>RNK]_:a<1IWLQA)g;[GYf
M/U>]6NK5@UI9Z#Q3ZM^\R\3c(@edC]PB:HW0F&62TE;[N/P7G(>&N^[D:Od6A5H
_LDXMM[Z_[)&+b@?BAUS>V2V#Y4X>G^7^I5>S7:QF4.[>E/E1YTgAeR7\GeRWEUE
&KG_HQ1.A_X)>F6UX^fZDH59<(b:Sd+=1afH9abQ>8EE21\;FG=Z#V@fY^PPQU]e
99X_La_7D#\QE-@5dHV/9Kg\556TgSML/AT45eCXb]]FV>G&^0^DG-QBXZ]G?8TT
7Y-8W1VaWfM]ST2B6Q/JG;SR:>7EAEM<WG[\a#89_DD1/R^>V4DbZUJd[=.Gd;GS
VbY?C>(EO67UZ/:7(/22N=3B<N8NT^b]82Y;LNRM2(@eYT2g[AL/2J3gX?1._WAT
MGA>K7O]97Z5W218(46a->Ba_2(:eZZVF35eR-bdLQ9WT>eIR406a5F;J8JZ]a_+
+H5Jgc:9/^3P=[<8IXF+A(L24ER]@+/]4[@AKWU?(e9KdDWgZcebGOdOTKdIQQRS
(--)___AZ&b^Bf?27<ed<f^;KHG5K2d<;?g?9/AA>JCU+BJ5H4fF:S_@KJa-R[WE
GR1]4fIA;FS&-YF_KPL9Xc^eSEG(]YCE&E2.]_-63NaNX<KD?DP0ZFJ2[AZ<_PdV
H2L#X-J3CG)BU0NLCW0b71_//2+f;[[b^Q:Sc_1-O-UBOK@f(]a,;N=+TF)/0aU1
d[U^B1I)C#BR05g;GL>7b=5K^S_EPf5G8.;M6KA:E],GgAB[]a)_R+/FA&eH/2fI
0.TX-fRD]F;6&=57+aAdZZ7:M6L+Gf&RXE2.<A-T-M(I:<C<GHb3ddHW[PWXc#Zc
d5A70=F#T,H2>SMV+F6>]EaP(c?J7;Eg+F+.@K58SA8]?f;[0GJ<.,-+BZF#f]+&
WUd^0.f07)O;d/@<e?#)\a?EHX@&V[EI<EMGG[3TK9:-1J[Fd=II4^SC+.f=gL)1
A0>(>/\C5/adDf1EA4S/(G2^.(T?18#68H\W6R\W7U-<(V-SOAb<WUJO08T2A7D)
(KJJQH5=Dgb&8L#)-\KH:CGB@R7?6UA2E,[W_0a2EL1)EJf#80OY,8NIZ@>,6R&8
b4(Z9-T+W@3F_>G^,cWU#Q/A88[OIS#JQ#09;I.=Z)BdAX:.Z?7#?<^X6.ME2S23
:Q(S8+.XHY^Y4;P1WF08]S,fH^PN_BFS+X14[fGZcNQHJ-=f+DD(&5)_^EKAZK<M
TDN[7+ffb^UOaT5]fQfG@T7P17.A;:7E]WX@V,E;<Xd2.UE#_J6#R7WBMX-1Ab^(
/2C9,H.GI32_30^.--<SLN:]b4aOJ\H\3,S7#1WX\X(d=(8L274AL^P>:U^#@ZY#
,=,N1UL5]Q+<dM_aSQS9;#Y&0fI@a4gJ7KX4.]><^JL@,.IAX,ReDLY\AZ5\ZZ+?
M@@VZE(_SOWG&4D)A4]I7W:=bVH6ACVSEH]eI8263V4(AEQDCHZRaG-NDCMB<0gZ
;>+N<6F?D+;WXI8WJ,=B#(<&//SFEEMG?(N5D4,XJAKMAeV7LO,Y=ESc>E?;#fJQ
?(+T;^<H_3ZY_Z9QGc\\5,3575f1cS/R_](.A1T#O)8^\<:5PeH;4eD4-1WU];#/
K[8->N;]5fT[_-\+)TZ;&TZ4c-VGGPb-R-]TX,SI_-?Z<NOfQKEC>#Q1UgYQgH0?
U@>+&FI[QK)E6R,g=Z/6YRIN-C\bQ1<d5CU__AW0La+=[[S7AO7UF?NAcNd,_^_V
JP^9a9HRVNF9>9d+XG=V0YZ&f(=YVBc:EQMR-Ce-bRC05@4VP=GDD[-92<F[ab/H
VNZ#W1.R@U^7JcdQf1^ZS]7I=b0b&&3ZN4MRD:]?3U[@Z+XA1FNRg#BAMafe+:82
Z>f,7@RcKXG+F\/NCRAWD4T)J=K2G7),/NO#M0@@H2P0F-KU7>VMB?A^5bCNeaKD
L[I#0_NRR]I>2-/:GTg&AUf?Q#EM?cAR>cLMdgE6H5K;3YUeeSZ^>C8PC5=RB_Zc
RC8?[,/:Ye[#RA7<&Be1cGY:_2]I&L_WITU<5@7Oag5Ef2_)UG&A/3P(bA,O+^DG
e)9f-(dOBEb?X/7Te]L3V[.1].Le5STQfUYLIJUgb8Ige0PD]>:W0)G^RK-\Q9#(
K;EfDUJQT2AH=ADQ[[W.dce[Ng3#ZUH1T[G)?F?1Y<T.5N?S.ELS4?;:O,_F2@2M
O>##P;W15NWg-)#4[DH/dWFHE<>)@1R]::/M1NY;FSFB,A;?E<)^^;N3S@@,?SOH
<8]-<V)XRLSY=)7[0/cU[_2#M?0&I)Z<R>0.L&,:U;)GH6eZOKG]6c/X4J:5:_>T
+cY<bcG)K(\6J9SE8@\cd#<EQ6ZOQM4(BF:dY?A(RRdYeZTV<286P1Mb@&BaLbHE
32X&_^MS_3[f;SNdU<^&Jd@+Z1ePA2W-+WU?1V#36ZPbed2G_SB[X#[Y+g>ZA<Yc
5NMV?1cX<2+,6L&T6EG95J?=<3aN__D<8^^@FFe;EYAHO#<?P]YW,2[M/9C.eH+_
WNH7X+,2TMUBLD@E5\b\:CeENHSTd_bTb6==RG>;/W(cA3Dab\[@YS^U=SHg9&])
J(DeN#T\W0)K1C8_VR7V@?fV].FNQ2Q?R@+c]fUFRX1GWY&;I?S(0&QND.4b=]\_
a^Q+K8b)MK3]]V5GB#F]ZOY4fDEV[T.?g68.3f\7YI-_HAGKYGf;dQP4?#?D\?;[
UfRB?Yb-SEGRXS]#WVHGB_Dg&PW64W?0+7W.Z?#3O\)I,V.K=b31?VZ8<QI.Jc8K
e2C_eD#9\&1H[a8ESQDU(FG>e@V^/NMTD7.;/U6G?RO,dF)5IQ,e+EgQ4Z^Y;A/e
\4]PU.@)G<9D0U5_;Fbf/a+ddN?;1([[GQ9-LV.Jd-)@f9M31E,cC/TK1O;BGLPf
/b:OdaC\Ze]/:.XdANdP#RV78@4IKAP].NVR5;0#/Fca5A0g:[F=aH,]\QB1W-SG
7C&8G2(YZZ5MF8f>_<=@47:NLLYY&gA3L(25:g1\Y1\K)Pc>N+32Pf@4e/\cF+eJ
e>_5F8T7N06.^1e0b8Bcad>+447Ra4BGWBDVA:F,:]fN):aQ=_K6-MA#,UY0dMP8
_=77JcC_J0HX8.Ye0Q-L3M)M+EO\(?Tc=[QU>##a+:S)20@/I53_J:&ZQR-6#H@R
[cS4)a4?_&/#DP(([KS9H9<X1Z>da39eBPFSN4MK48UfGa^,VT\Q;eB9=eSTA2gI
(-5L@/TNaW.fFKBA+&D=TPQg2L\+\;>6UE^+g(S=GD?NVT1Ta-VT6:4-+AO-(d8Y
;V:gL87AGNS1;R6Vg6>-/]a^,Rb&=F4M_I3Q9Ke8&9e1K,R0WME7KM6L<M).cTM6
CLE>Z#@(8g[GR+ARQSX\&B+:FfHa_L.Z?+C2AP3NbY8,gW:LIBLI@)N+HD,L-+[/
f9_/I\:2[7Je#AK;aR-Y@(HHXPAM@OB4)>R#2d2[6cP;N1VUMS/>0H=<Ke^Y0aEe
OJR:03E.e4;G8L.:?^J5<Gg8eA35&=ZEa0Q>QGdg3PP:5ZT(ZKL=dBdF6K])(H<\
ID=g=fY/</B0I:TKW;()]8bUWFJ8^]?\1N0-UAf.I]f+TaV&L>(Q]?+95_baHZ?,
N87Y&8ScTc0@-&AZ6.)YI3X4E5OcRMOR5RM/cTe+50G=(39K/[R)45(QM^R[JH+5
.N_@(-1HQ,#1\K\X^Z\ZMULW1\:QF+gTU2R/K?>/VS5.g,CM\HXSB5(aA,CSC6[?
^>a?<J=O@c1?K+W#QRVIRVAS:H8\Gg72Q(]BgF4U7Z/Dg?]=;8#.6YYH,dA2#cKH
H(f7]UQUc[#g1gARcEbU)0EdM;eZ(=3IaQ9>e:9@X\X(X7QE,Ig@:J:X]P=3OUP&
\C.B-3GaL/R_2(.Kc)ZA15U9FCAf@B>1=#ZZ=Gb)EcC]>a75J)1E,UcFA\6/X13-
X@0eK?g-#B_NK.56?DG7L:J.d3)P(W^^@E7dJ=JE;;#@JV#1++<^MdgZ<UPU?Ibf
_NMSMH[Y//bBb(KGDG[[Zb=GCaJECVK#=Tfc[@Mf6[JB4/8V_-T3#@bg8UW;C#++
WI;B2e(F?;g/A]E>(7R0<>Q(e1.(OR=BdWI@Q[LAZ]Q8&>>ZO+cQVXN+/Y@a8gaX
^=:T4\0UYOf6D15c9=AFV/NFdAMX\,)V^f?e_OP?4K;adK&c0+4<6O_cGY-)UfQX
X:0gHdBX@QgEH;)@8)c8#IB.O-F&Y]I9eK6Gf,2;[W8I2>2=M(56UJ7D)PZ@FV5]
eLEON,)0][0]=7_fG]DC^AF)J8N6ZKJa(F#@,6AFK?X;40;MT&YVRT2&eOSCBY>G
9f4MZ4cdBf4eKc+.Q)_Pe>MNRDEY[8X4J+TaCag896M##Y)1U\0bR=6Z2c\bK,]8
6G22]&BLU>DJ+]8TX?+E_:R.&9/P+Z--JQ=G>MN2:9Gc#,eZU-KUY;ScQ709Q381
:VE@ENddD)P-7gd;:U&JEY=EQdRI+KQR4IV<,@Reg3S3[4G>KC?HO6CcQ&A+9BKX
VKV\\D.-PU9A[=36/P@g>I=f3cT1A[&=[IIZ3(;CQeS^@D=/C))+EW<=#f9ZMKW&
+?]P::#YK#:]JHO??FPRW(8&T-)\0gDYJ2B]1Xf@Sg.VLeOG_7_4@_W:881-L+bc
4NZD_MAR4I^abY/cX>6bYA4(>W=J_6gMd^^0>5A+X8ATFD727X462@gZTVO)E)+V
-dIM0J66IIZZ[R8HDcB53d5+1HS)6)6a:g&I_D/U_EcZc_4:@?YGV;7)JDRO]fH7
G1aPXY/=:(T5d_LIWTNTW,YKKE^Z01Da;0Z<?XPH>XXQH?[\+_Pe7SOTMfX>=Ja4
U=DM,T=<TE;09WA532L<1>.8#MD83,H?fA+,4e8/V@>C8IdY2-)37^7fd^;Jb5?9
eT>dNKO,]T>aOG1Ra+W+#W8M1RF)DeG6(3JI4=UY)GfE-d,DL<[#9Z+1GbB,)Q>Y
B;]O]dLKO.PS^W8-8T+38WNK+,MeF.RDd,S_agK3@dH^MbUVJaScg_GM_XgES-7:
C,RV)D6KD?_)0S;W5^^K5d:\HU\S[1A.86cYQ72.LD<7(ER;EDO,-BdT-@LV[M;3
>bbbF[Lg\)G+.0d#6OREd@6S(H\#+6Jg6#2Z.GR_^2-UCI^1R80MQ2YS#><UBOLD
U79VIH44/a7P^V&&M66ZLb3B80@&[Q4Z[S^6YOaI+#b^M[bH/7bQ3S]#A:faZ6/_
?2e8L1Q<,d03>[;FQAGI)F)>?AG/>D#X?K#DbSOYgXd0d-2I<2D1A/)JAA<1/A8,
4;6UP8-IU,WD?3/R@VFP99=+K]X5Tcc:K^K3Q(<#MYKX7L\37\J[0(OPfSId9_F;
LWT&f(VeA9aKdS0_:H\MEFH8?EP)g0>(,eQ@BVTd3]\UH4)?fZZ,7PKB[gaZ#.a3
JT<.aH-TE#7:^S9#>f+E@_d>=34aAY3Ub[?gT>N\]EMZ:Pg1864J^I2@d2VB3Cb1
f^3^a=SL(21(QQ&@URbVcg;O.d]4LUM)#YY=M+0/P_]W#[)CY^:H(MH8C-gLQ)LQ
<R,1]M;5M/BBL&;@U5X0ORU.SYM:4+F):_N1#87V\@5I&K7?gEJ8a1ZQ-STd22YC
&;dEg[\BGKO-)ARQG9-a\P9O9MD)5+f-D[P.AX\Ca/be9c7f,5Y#)EJ?7gQfO([J
6U&T-T</&/-)+Y<-8XR8(E@9L@CHEbE2AC8X:(-I,6bR)YQ39[HS].OPWZfeHOc=
28-PMUK\-G;-_/S73RD@fCY72[,9L(&B==&EN&IQD11@;UZ:-Q.aX^g<S;B_[BXN
-1=ALG.FTc\F#c19RJH>&_#P;YN5IL+TRPQccEN_7HS/HK><D1<):DEdJ2OJWVSa
g/+Da&b9PS-YNA@;aNZN]&=5Uc;^3(76Y)0_VQg6:^:d_0f&XSIe7.LJ[IUfda/1
F8K4FY)59SQ3T[QF2UbRMaUZ=J&3c#JON.-W/WPT>W.<7Q/RCC5T8I+)H^Q9Z-=:
V(U,/6=X>@,a/dM=TG39EFZ@(N_dUGX9_N7Y,fH)@):,fW;0X)XAKQ,W[\TMVaC#
:?W_e?.T=,<JHEc)c-DHWbJa0QecZ.MaP?MJ59,7cK_<1C1RFUZdKR=T\.@\[De0
HIOZ]F?I[9IE),7J6Og_]R0T2TK+[\#F:OSPS>(J_HTA[NI8XZEe7#?eU6WML@UN
5\J_FTZ)6?C3SF:A6_NG/P-F3]\VZ^,0/NfCGH^/S56+@8JT@9LVX-.Q2Ag3R7O<
b=ZY.D^DFQf+M],aVeb8[(@I\GQ9DHWX7bf&R=KYF&I5)W;Q_IVIAL1K^^E<_-gE
OY+HT>BM5=O;)b6GZ86..ZV<.S;UZ5O4b<3&VWH3,N)7b:P;@9REeV/0_cR=BA::
]XES5cJeCY-NH:]c^L6&39Z[EJRYLW[DI0d,c,[9>95P)1.#8AVLRgUSGW8ZRNK=
3EUKHT?:>#F,5)5:?LCI.B[>6eKM3V?4_Z&X9=_YJb4>((UJ>@SU8D3Z6OZ2c[N5
9FBF]9B^_ea?,NO3=,M/L)P=QHa(&N&Q2>QFdS>UC3::f8;:\Y-faf(d87+59H4F
:7B#G#IM(a5JA-@+XKcb+JQ>]LY3?f]Pc0FB??^_KE\IW\D]fMNH50XL/)FK3N97
G&\5<9dC81@,74_:NcJC?VXK6aR/=A90a>#=T.:@RJ^G:3+a[=89N+PEg?cg9Z#N
Ib+Jc8[./#aeRA-_N5YSOe,+N#[Ca/UfcV)b#bT7XMKAQaAAF2LLF8@0+DFbG,9H
B5\1ZY(Fd@/X3O9+&@1REEEg7P\2P=&[6/9(DKCcA(;MM7Ze7NXFI+31(gJ(7R0A
D=ZX,.[>JUU\_YIB(Y\,8-G#XN[)2G.X=a-LJ]LIXZ@aXeO<E+_CTF.8USc9R),V
9<T+eQ/4^4;I&f7?O4EFaBB&g8C9\H/8?G\LcP]S\\Uc4fbE3/U&82/Ta79??JD&
2Cc?<M-K+XGPb/IMPKAFL>)])_BA[e:X;Da,#E:e9#TVX@gS7EQ1)9c7g;N>EV7\
J65<aL;;S5=[g)DMBZMK:OEP67>^D,;geOZ(9d564ZYdFV=A]B;#dB#9_KRd0ec8
CEcZNYUR&cW#deJLG1#[\8Q>23da?I&@Td,OO,0\J(Sg096].NHH,KW#2#-7?FO^
/]155gb84<N=c6#L54V?84&/R2BQ,-=LCcZNS?D-aa28Q,=)^W&4-L;FWILN70Q\
HFCcXF@,EZ5eS^]KW=]7,=7bKV3STNc6T=\IgKJd]MQHRI4)U&^f63).@+&)=G73
HDc]1J=e?NeIEX\&-CM0@1QRK)@dFYIG><8c2&?IF>L2c?C:?3FfM>0W?RaR-5A@
>TI5Y@LVeg&R,HgO_[5V_[[6MbAGPOT.^W0BO0CD;^NL2^C6aIHS)<K.P21fb86<
\?DPbL0Z6N]:I_4WUd)6A?QW1Z0Ka9\:BKD63<#?>_;S?SG>6>X4Z6(<JAG:07P5
Ie;EPLDKYg>U-+N8/Z7OD\>a)R):))X.GbURJ(5?EXF[]XAM:cLCd4R/-?:V9]_f
Sf)J[)]EM8S0.(3^\_?;SQ69+1EJJ>R5EP?KLUfNSQN]KW3R#fgJOc(3A^K(I>--
KfPJ)?&T,:)bWM#Zc&>@CfMHK^OcJXBOdBY+FF)eDWfLW.+\ZCME#-5B(;O;_Cf;
X:?P_N]H2dC8Gcg,e-8a^c,SX(SC(DXF+IJ5(b]d2#b<L?H&YS6g4g9e^4c&g.V_
J\0[:8+(]9V#<0MgM)TD)g&FD(0MgXF)#3g5.0YBU@M7V=V10]>Jc?OWPR2A.]5D
[0D>O4I.31/,abU>B]5DJ(U-S];Q+E=<HN2#H:SGbKW_M(DM^B4_MW_fEM9G33Hf
fESZ,8O0=&ADX:QfA:O>CMY/(b,OAO=B&#-c\Yf2PQNV\G>7TCd=#][<NTFa#-c<
-BR_?OS_E=Jg,.dEL]c?9])/-B?D<^O,SP52)XF8,\C^L,BG7,M3K?Y-:Y##K5X_
TRY,IS;?ZTUUE.,)cB7)ZME/.I?+PWG/N/8bG<2KEXff03HHD](EbJ;)J/(Mc:dd
:_@LV87^X>GN[_^T)3=Q)GB&#8ET4AY&?0J&WF[;7[VV\H)XRAST)Q+EWO=6C&EG
4UJQN2LZMME1d>/B4[2SJI/SIA_YM5aPeU<c(cSX5aEX_FNCMY2We7#[?N+HW9>:
<=G?K+MXPW/:W@0I6D))e=4T/UWX,?I8C+8D?2(93(L4).ZW(ROTDG/ML+.Q:R,H
3f_>:[_0S/BFVMeg::\e)Z3;&9#6I-;-^;ZWBMB?6VXUZ[ffWAI[dA\=-U6&TK<5
HXW)^CUSfG4cV>\9FZ6_5c?>FFY@YV.41a\aaXF,BZ<GC:bg>9-2]O_/J>>R7_5)
I7XVgFQc9aeT:6)cRTNN.Fed>627T1cXCL:3Z;1d;g0S_67VYU#_?a1NI<YWe9<-
ZMX9bO?8Q>XUV]Z?<Q7XHO?7\3YH]C_^7fU9fR8[V<IfC#P]c=@-@:8AfE6B2(LS
;I8?F745NGJQ)39]6>?FB\XMd.JOdZ.@a1AKA/]Sf:ZVHAQ2KVaWUTccR?&O].L@
1@,Eb8MY;;&C/dDT^U]Pa020+eZLXK1S1+,0cEA:/@N4W[g^BXQ##cJ,@]5XL?ZA
.\L&21[^52O#gV8H:1#SPaMZHY7&d9@L2/N\a9:^MHQ#&&:6M>6C)-XG,YJ3(E)F
c<=&]S/N(P6KKX=GW_ULT_FR-],C6gRf81\5.Q01&,#B>,@GS81)[JYLN2NRK>(7
1X:.BW/+^,QFD:TL&/f0>fPRbOC@,@b@^c8Z:YaGWD/^QHZdMPCeQKK..eAL33VM
&P:KY^a>ZNW63[,6>MFfbZO7_(;7_G&I9aOAXY=BU0EXYDUV>,>>IAeEKHP_9O9L
\]gWCRLJGA7^SUf1bXZC:Y(YBX0+(Tf8e,&D,UL3.LHe9^:-:Q1TbNMegNWPaJ8(
:O9+1##Tf/H:UN]3Fe#:5S=(8<?]N)f;&2]F/\UV@S,ePM6QMHC3AZ#KFe77#,R1
+VTBC7R&g_TJOY#Q>fR_JQHUS(WO2T;:WeV0fI-cX+;V/JN>TDJ7>G6PN0DO_\aQ
/9fU2@(>/d[5PV2[0d#.RfLS].Q3F)Ne@;<9g,=YGM;O2M-^+R##)?_b6IL#G6MK
L64ZgD&[]S:bXE6_e:fQNW5Ia/)1N>+2=D]^H-&@6[WW:4@DE8,E3SJF3[G]C2L2
@4e[B-AH-=_;@3IG+cg<>Hg>3.H/(UD&]8dQF_:X,65@Nf1(Ad<L#:?F.D8C^)W:
\C?ORVQ0>&2VPO#=4<+aX@^J6\#RQ2);dRF]EYE.;g7_D,]c+;NW@1JN\[0Z@T],
G=0QR022)XLJ:bQIH6)QK+b25d\?XBXRN^G9ZS1CZH:@.GMHScd@XZf@^>JI+/gS
-W?HEOTgbX\;N/b&GQbXTNS+ELFBB-5,7a4F>)64W=Z;+bZIgXC#?[MLP==4F3EY
\d\_A;P<aY7XS/#Y^Reb^cf/(MXQ;Q<0dRMDb_ZN7@9\U;9Tf5ULEB_K+2:dH/bE
/0LK,g.=Z5b-eOTF]AF+:0-NOUFfRHKHKgZ,AJ2C,ZNK3c22g)eBa^V8[0J\PgKY
03_CWcA]]A^B<R#4?M@710H5O5eL#-O;-&[-[M>TM)=8T;=Y:e_KKIUHEgIY_0)Q
[eXCQE-]=XH[3+X3T18VU6YRB>^dHC1].PZQc=TLW4K&Uf.=F]Ge+[X:aV/IdJR9
4<9]KK.Ic)6g,9fF8PXOd0;W9GSN4-9O5<]@J^Q<GMN5D\,NX0S7Y7IT#0N;)@KU
/@1#C@M;.QF-TTEgO8Z@7)0bScC0R5fa[,Z++8.?L;?Q>TW;YV),4KIJ#AL/0+CP
+1#G3)@_6dYFF7>5N4-g\TU.HQ=bY_=I4WEU]F5feN4D4[4=>0:1:dAW80)OBGU3
KeXQN;_8F^/Y&91D<M)O&E\2<Ncg4LU3-aI56-f,:PK[EW&b6.?QRJeaKYG.PD@K
&23cec;O)C)-78L9VH\:g/-WR4DISS_3J;a67g]X)==LW06;:>9HHfN=2(Xf0^7<
KBdNA^KV7;FS&Je+da/.LQ<-OGMYH9@aPbS98&28Q@e8M:0MN9O:#XCUV)N_-/)C
FIc0\b1E0M0f:]Z\WRg1:V)R4\UZ:Bbd7CA</N,3+?Z;dQ@VC,gMFRNE;O40S(9\
#&dX:.&JY12ODS:??@<A)/T3JJa;9@4>^H37AMYb5c(8Q-.dYLO^7a=b&MAAc_2U
<&]A<TDS:4Ib_U=@0\ScA<R6G&[L-L&d[d^N?2?@>.=(@gaT,g@d6Z&]Y@VdfOKL
&;VgE>K+AeeHLJ(f]B15DN0.I8J\UMf697IdQ89=4/Ha+W/C+[1146Q7_V;C\Tg>
MNB-CN3O.+f;UG\V^NNG9ef^@+A]G1Fe=bY78Y]5CE2:bS_BU/F9UfB1(0\GY9<@
2]LgH<6L?=(SS#0d0L4=#;g](MFT/-2(aR^RdF121=3U>PXH1K#941KC^@B2#=OA
U:@J-eNf8>SJ@U6W2H.B<?a(dAg@&V=^Ba&@QCSS)U[f/g)bC;b2DM]5>CPO,,?>
XBVd#W:=Gg;B47\a_E+F1\bg[&R<X&GVb/0aP4^FTVFgbLM5dDf751#D1N3=BS#6
0Q56^(;3&3:KJ#,8:\bSeg<0S6INQ.bg<1R>-_ed^XX+H,L1):CXD2f_>MXNFL#\
6DJ.2Z6V97MM5_#7AE@-CNEX1_TKXOFe_#1#GSCWGAD0SS]86J?,>(?[OURP06LY
TL_WZ&O(>3_b.U7HMW)PLLUVf_?WG0J2gbIXY5Z(E6dGCNAG60O>a[SF#24+@A9I
WLM7b5BQ7ARU<15fDL&5=F(F2cW.3d)f2EA_b2dHP)==/>&ZbG3=\d2R=[64#a.J
X4#[b63X#@690.-)(^X:=D;+U\2[0d(]?QZD@>JgT)SR0G1K4=NV8Q..H;e)/0.:
0ZH@aIJY).][P1,b/&K/ZQDFHf>R6)2Z+VN5-KDXG3P(T51<82T&(?)U?]K;ZL>I
3I.5B0G,G_\;C/3WI/25MF\O-I5L,Ya(K=1:@IXM@-a(M.gF8C?NA2QXMFgR1>9Z
3[^R,H@9.F.:b9AM.I)H_L?=1^+NcLKb/T\-CNK0;(1B[d==b2X_[:AK]Y0H3Y)_
UAR,WH1^#&M]O8fHLa8&+:&)6[=N/L33RH/\<+>I23\LL\W=2ZN&23/3,@ARd^Z,
<DdP>e9LET+X9?)K5fbN.>P(V=WRM4PBE>8AUJH&F6:4Z2LbD<WfS<Pa/1[bK7Ug
fW[-2Z.RQHX&F:8Ae2:[B]=A874SMRLUQ5P,R780gQ=Z7O80g=CC+3XZBY,HUe^L
/S3B5U\28&4QJRO7\1Y-F7?aa:^&VfO4:B3U00MXD(5.D1FN&1063KAEc0#b^+If
Z8aW\,7I=C_+]Sf)^S0_5=B533aL5KDXOZ2OS2/J\NL#OQ/2]8VN<F-DcK,;>+)#
d4ERLI7c8M(RIS_WQ?gR97U0+=aONA@FLS__-XdIf+(.O.ZLbX+052[cgXJT^g1?
+WNFbV8151/\P7L.>^A,.SZgcFS:g8aFTBZK.MIHg;\FAUYg6<ceIEcX/CU^QJdW
B9L57eA]/.WK98cP8MYa8HWTd]Y(gg7&4MO4)TCJ7>6gU@1I[(dK2BPO\-SXK8,b
TcR0Y]M_2@>1:^-MGPX8QX3TO_6EReYQ2LAS/HWdYX]ES]b[I[eD_VO,9I9H3/Te
>5+#UL[T9AQ\Q1dPD+@?<YfO,-]?I94PH(N3?X717@;\T0__cM2:e(W2?gK6::?S
^?]/#^8>L4W^Y,Y7Ddb:-<>KP\FL:\@C93QFcM=1C54AGf.Q81RFZ@Y[]6AJF3_S
LDUG_;\c#SCUTb8bgJe4473F;ER7gD+Uf)W/dR6e:DG3E_@A5(8ULWN1UXe\)I>.
EJFDCH_XCRK,/ITSI__R:EC3^ZeKNg:-M+.JY_J<F22A;]+8UUfebN6#a1,I/:LL
4N2FBadIS:=];RPCW>,7db;;?PW\_&1/<^105eFN=eX<[#FT)LcL]VII8QETHb8T
61K;)&??[R?#Z68?GM4=]P5C2/X;aRU+bTPc3&YN8A(@aSa[)JSbGH1>c)66;.N[
T4\43/>EIcNfK)P2&LMK.[1W.=/2HN_QF-Na7,:25UNaZ#KKFU&&A33]-UAJFM76
Q&U/]88X\0&LePR,;W@Y\Nc@/eUC30Fe[+Ne,H+D8T]Gc.?@WJdTW5)ZK\UDLI>_
F,0&5(.eATCSBb-F,ebW]+bgRec?f@M:>c:XIW3)bf;GBJO2]J#+ERYTYY_:(Ya1
S?_aA5WF:867&&LdF(a>B]/,4]CA3.UT0XF0TeVJE+Ld2;b5SW[+[DU&b8ASCcZX
?X=;8b9RYeOaVS/0\C6g4\K7/9W2&(5(LaK8-Z-2g>;?c;)P[^a-O<WK:>OWLg.-
H>ZP\gBB+@>]IAJ(#f8a=M\;=7>GVSe2W<CeCDf1YFB9Q&gXCN9SZ,gZM3M1+,+Z
<M8d&T?\4^@/XQ\aASUeRB6LU:3,O:5U)]Q[a\:Q2eX>WbM-\-?LJ4AFSF8(9D\@
FET7g)73UZD\MA\Q).<G/>M=V.I)4LWW_HR-]VfXUf/HZTN0\M.&4f4XYYAB?(5N
56?-^T8XL.Aag,AZ4>:U<S#JagPI:)EW#>WJMg]DCS;7T/DW>c0Q#T4C?6D6]XZY
MWf1&F&T6f\2f3HI9g_+Wd=E//d?6+bER<BZ80N#73R_;A=V\#-QFIJ0.-\@6A)\
>?OG@QXHB+DScX6L5F=R+:K&89RVa@:&3:F(88W=Vdg1[N2AZ:/@\#4S-Q2DSUV5
IeA9#UW.,M-1X/));ALa]#875H.K&fSL_23691OLYg:XXD7[(U?6I5UD/\YKa.I,
_0^dH[F<6[J/WeJHC.O[XX=ff?D^>1+#;8b1.4\.H;U[+)?e\6@\dL6H2QWK]=Q]
N52-]8M.OS^H[W[=NUQ4K3D[4N>KWc=AE1E9De35;eC9T#S4;NJ9:\IBbX;_YAF=
Q1D<VDZ>Zf4.=M@=VU\1N&H17U]Ka;5_28.IBKO0e_KE-I>UU^.8KC.ZWQW;d/X;
/HC:(LZW=&\CE5^(b3/J^g-7BZT](0>b[LK8@\a>Q2L)7REW]DHJAa;BY:AB,N5I
0e#f[^;F+E->W;.7KWAU,.8MdRW^X02IZ0@=gU>3[3E;S2>9PO4QL<@WO>F8F2:0
KeFFYgdU+R^D_BE-C,BGCY+M<f96#CLV/B->?;)J-#5>8]#KPOP(<87Z[@eC5=S<
,JQ<&:B)&QPI:e.619+@H\VG)7Rfb2>A#cND>c>>FHa=^gQ^CMV>IaN73>E+\Yd^
U8:JHJ4(-?<6dfKTIDg7)S9\39Ve,ZJ,??Ke;J?KYPQDA31.3?[bf;M9Y&-1IY@D
X8O:>0;__4cC_3\-bTTe,2U(+]cHDA[QC>E5:XA/eK=6/DRd)8(S<LGWFO=#WZ_9
Y\N0Ka\<^2cE_B1dX\9e;[4#_=ffeWAO2NA9T]fLK60GPf\+G;gS:H^<\2SYO56F
0X^+9(2SJ7A:aX2D:TI>>GBDFPKfcXMB1QPPQHZ1&CaQ/L_f]7MVXQ)#\^[P5?Zd
))2BACdaS1B\eLQ]-U\MY:>=b]B01>1^\DB_7B0PS3cGg,Pc?IV)3BO/\;O,?bZE
T?9<3O]:R,5Z-J(d@9B3&978e^c7Z<NfFg0D#R/:)GJD1<=Y>ZJVO-2G@0L1]N&5
VVFXVD6?3?3T6HT(TE7^:6AP+^3Daf@,(D93ZM,?Yc(gM(2C32;-^cQ6eC-d.7/5
<2<K;aCb&5Z/J\QH]/2CIeg5?=:^4=>QfPG8e-b9Q+FB)Z+1U^[6G([(,&+]4-K,
W=7\;7GN<7Y:,R.=8cbO^1VBM<T:J30(NG7AO)SQ[(TWPJDK+f.4Q&J^E>V528C,
deU<GJ-Z,V.?^e)XJ.:D,S[N<R3e.gX.;U7<FB\WL.gFV4->gH(A1b@<//UUGL=1
f))C>JO9VA9=Lc6U<4YEFQ1K#a+8V64]QcX@[63)Q[W2BTI(+PB-)<W/L9J=;BN\
]D+DaXfc6M&8bO]_&ZINW#1d\P_ReX?BU+;UbOL5G&>K?1++2-AYX4H=E);Kc;=]
4G(>+\HN1=[\,[F0:SY:.(_gHH&Bc@V5R9WYI@fa+&/UFO?:5;R<.<&G+)^f5b1V
-d#X5BY,]78;113#W926B/+V(K3.97IKU\?F^&_OW2,@<WeeNRN0QC?WXMN,ac8L
:3LX@<SA[_SXPDBWXI@Bb&P3O2+Mf94_N\Q3\VTX9@[)[NUG]5b.Vd)SE?HTF)8#
\,d7Se2ED]).aN64?##\&B0Ob.,cDdSQX5RA4_EVO5IIa[NP0S_<2H6\Q6]XQ+eO
#:]0V,6caWAF96=JELOQf6=^0;#W16H9U-;C9)aef7)XGSNO)2YD;;J8.XW=.YUb
;YH<EX7A^^))R:;=^Ia=L+SOL@AZ?Gd4XIg2PJaAZA,:3/O[3,fL)L;g2HY-_2>>
Ag(KVNB=+5,XgA(T\PNe^Y^P?4S;dJY-_L8b)T\?L_UT2f3f(D1CCCQJ>E<?PcOP
SKP]U5=7JQ>GdfY;a(SF&E2CNg=;0K1BT]9[d/QVfBLS\5O&R)VB<]f#Cg>]f\?&
@A7[RgK-+^C.IC#6:TI-AeA>T]X;EY9T)IDCI59RI5=d95,9W+B=KOFZ:YRN>&=8
eVSc,^?bR\J2bU1c.@U_+fg@73EJeLA.IB<A:fI7:>4fbHLgBF\V[.T[-&QA?c/E
Y6a]1KWK,.<-E:NYDeebQ\a@;IZA)UKF\MH&+&=d5#K-QCc?)AVdaBb.<cdbTUDF
WQG_->@>eZ?(Ed/NHda3b,Z#WKHc5O51)KN)V3@:)R6N[&FSZTDCPPMF>\:)OE3E
0=7_NVA/QeTKD2?Z=W6T<4>5fd5/KJ,_>Q+_\=HG@JL[F@_&K(#U]\7K:S>HY_56
I_,Vb&Z;I.DG>W@H0<O39ZD50LcB.9VDFD&V)d_-EbGScK&46IF^W]Y>G(6>gT1g
SJ8,Q_+eL:,)O9K)2eN4WBeN:+#/MM+&Z?/+X?J1#.U.fD47FA[WN03PY>2^X6/\
VLB^_@\GBESK58?#2NKf1E-F7,=YM5aEC\F;ge\BF+\b(2Lf/\]I#I@23T:B6f#X
EbdOc>eWc:W8DS)(B)GgZgENZBCC2)4\>Q4DMO0R0e1;RAWX[:_//]eCbb/gf^0O
Q3D+bgA[.R&L@D,:17@b(R)CAKF465;635HI?R#&4a:ZP;^2Ff#_6a-Ud5=7&[@P
g=E.U18^1VD>d44eOS/YY]8>=DX\J(aDWDD154abD&PbR.(V)EIJVGM-S<VEf5,X
^b-9E&H(JP-Nf)]N2F;?-7X6C2E;+Y3322IM(&+FI:fRBNG]V-/]bg?A44e>cJX_
+3G2a2IM2PWc(>WQAS\X\J>#=3eBO;c6bD/PF):(-b#;17T&>_X-30+7#a9W4-:L
0T_A+1M:V?-O138T-_=PE6c8K6<C+/=FeAUVZ/GfOV2HMQL8B1N&>P,:.U1L&DKd
EL4[P..d0F.Ff@D-1be;?;]QVF<F&B0ce/d/R&=IbG+a9cVgOX;;aa#15T3>F-41
^,bU=UZVaUK(?H=JZ-B(2N54:6;<b92MDURYJ=@K.X5_\AK&F#5\VbVcQHCFLJ.(
V5-(SM5@IUDWR3,gQXW2BP[9a&c(AgHXWVIYR\EZRO7LA)M4N&e+(:9+(Y?=U+Sg
U(G0C)6-,-N^-Y].M#G,Z=P3D^L:)9=e;OBgD)C#48/&L/QR(f>gYBI8)V8W1.Ac
I,a.^cX0/-3__ZdU46/9DbAf/6dS:=2YUe-d>cD;(\W3V^QMAA\aOPNac.RU^=VG
9db.9D97](g8Q#I96#A?LQIO=P?F&,:Y;4U:VUQ(4-:1#8OZ>/Uab]5bg#SAD6@C
?[XJ/0[^_DD1(MHH>^(^ebL@RMR5=L1<&0[FBJ_ZA7S][KQA&Y-HMKE6-N/.gR?U
eI,Xe0KB-PQP+Y3LL1>#L7.CK7#?<4R]RZ7Z0@;,4@.HU??(TT?a:&2V)AM&,KKZ
EG&M/P#aOUFSX</Z]ZT+AOM([3O^M3Y1)@/,EcSZ_4eJY.7YN/_5V:,3]RA4-#b0
N@R)>O>ScNNTAC/1d95RW)e^9-M(f&9,IYgTL&T+&PCX+[4;]XS557@I[fD)>^V>
b2MN0@RO?Xe4@b\LBCJ<-0CeB:MYcV8AN_NdBU=.ICT&cE#\.<O,&>BW;ZW0R]3/
MCZLKa#Q7F=e.M\+T/fG\EW_;FU?XHWI:-2b0BFCJ4+Zf[G?fQQE<867b5YT=J,E
.<(\X0/V(D4aL:)4<Z.?TH;1/GOf.BeP463dg/-b,,GH6c,+\+_gC?eC_5^D6H.A
[&],87b?c0?[<R/c[,0Y\<eREDC3Q>]d@O#?ODQ#Mba0&=E-U(UN+[)&2=]>13&7
7CB>MK<F1C7/\@Db:4&\K(YceCV\K3_0:AYTD0&5J&>]1U:)>2:E9,+YDIVL:[e4
6TOO^]/+[N]6gZ#c#;KWYA-B@e3(bc)g4<?dL[BA:(BI2G<4_1,4B:1f:b;f8dgB
XOPgHC]5(06WZ9;9RJTI/-O:/^<[)&\W-WEW(]9Cc2&CM/]&#G^?bOW^g<[L7LF/
4D^eD,[W9QecTY/16<255X0V0J_d5e1C5?(7MP4gLUaR\D#=Z:=E&+BPK1eY8^DW
eKE-S[g:FR&Mg8+3IY=&(Mab?D9D0BX>cgSKYMQXU:&fV7ReTB8Qd^T[6?7OC6DE
ZA.PKPFG0P-DXUQUe8DK(:LD^COZG-7FY78P-Y=b]8&L]\g+>BeI=SH_8@UB4DKN
_8+d6gYCPV2,9J93?MQ#6,3PL49cQN(Z=40)YG\cKR7>/Z-]Q<UN,536=;-4CgY=
2dR93YgWJdcNS<T.[(VR&AXO<bfcY&F)97LT-+f4FOg#WedHcY>eR4-Nd,W=_O][
KA^@FOGGNT(DOb=+bNbIB0024[1f14]GF7O+):CBdFgI@6d,B[U8a]Y1f0??W(X0
>K\F:VcW^&5OU>6e58,3(31\4PU:[Ef5QHR1;JeRSXRBDA[ZSB@[SfZE9RISLWLP
2cGdR_K]fg1f]MN7],H_<16c7P<WL_8(#CBAF+fNKa9F13M(?865+Sb?>5MM&O#2
.W)VT[HX74b5Vf9&]SVYgOU7TWTZ=AcAe2>^f>5L&+J,Z#296\#=gR0./&[;8]\G
_OHeN(K8PPFL)6)WT0Of;?:T.JBY:M:#WC2Og(/,IfRJ(.I0a)&c=NOgFTEK<bI,
Z1B-L-g<@)1/2b&D6(JF,cZCeGRIcWAHU><Z0[14JSY#gbbJT389-EI>+.G3DXHM
DGdYB&3R6Sc/83N^>C[M5)HGW<M+d8->0eKA(:aBGW\WYGK@:VNXR[]H\CgJ(L.c
1-Qf<bXf1P>H[5_RXQUNZJLGbF5N01D@P_K=-5^P37(RPf1RAHa0V@U;=H)cG(GP
f6@Y;S-96efR2][OJ0?YQ,aT5-Z((HOT(7OB:Z3I_O&)WY]Q;XWK9/)WND^:]0A8
Sc>1_,K,<X;8a?E?R_D=>3RVbbB/RGJdJ9e;EB>K>W^3+]/g-R<]aW[IUdf+\382
3CB4(+a]1bYL^238.ZdP981U5?Q:5=S&+c&MK\1XQ?;#(E_eL]]WU1#cGbKDYYV+
:+L4?;NJ0E&V=bEB,D:D;;N<7Ud-;6O/<.;]4U&_Hb1I81LLcTWg=+bA8P2eW03a
9[G/JFTQ[([\SYc=2<WRUCL-CF3YZRZC]JX?H5>=d]_]A:PDD\D4YLCYY;<eA/)M
GQ=V_L[B0R&5POJT;&de@QDdHM=SS:MI0AT]Pg<_?A1AE6YWW@_(8[1H(Yd8O;=T
fLV&GQ8X4I<&2UIKN8cK]6)\HK9>S65:Bg^G:NLC7U>cPY1H8W:1(61_K63VFDf=
>@LeP;^b6&/WeTf6\N45)L9^aW;aBAFeON#7GOI8.O(>XMFEJg<=L9fV@JX+.>=E
[YOYKW6cW>>W60#4-@L/G]YA5_ZET.\Z+)O<ROU3M_34dcV+WH/CJ61UWPMB5=HR
O-E-<P7/b(B#UZ-MR[X1]?+TPS^.PD?bf?g[8F.VL=&FHF0dLYBB/3UX<c?I)6?A
Gb]IZU(<<:86[=Z/)MG]K?U(M<APLJ3MP:.D,?-U)a?,5^6]G5_9S:X&X^SD#VM7
.I(67g/X8]M8&IS=5CP76/#,Dg<DG_]X<(J4HU5WKN7SEOU,61>-AH\c]V)Pg;J]
:,L-GCJM,e(7@/3D1g@^QH(g=@Lb=Cg.XYa)630;TQJX/I:G,-W.:,>F^dWeYW+8
=QTK43C:@E&c:6)E5BcQIX)<89ae_d/&/VWG/L^#10]TEa:@LaDSI0RD\#dbZb]>
_,:1U:CVU\ad,5Q)@YU\4Y.a6:=SI+EMc)JW5OEf;Q-1-dDVRC6d4X=[8#]GN5UM
B\QYIBE(DD]HfCeDP?7>8VYNCN]JCNU67-<Z3gMGN\2aO^LNa-\)4476_g:M8Y\,
+.??SfR1WO<GLQD(\56.>:c,B5,0+ZAO0/LY+ge+3AR03[eOf-gD]KBM;566b5\6
7CKK?aGcL2\?NI]7c(BL4<9-(NPL51\IGT>81ZC)AU5OLC9[aFc&S<If4^1Va7ba
J6<(5<X<D(X4L#2XcH:fCDZVX:b[I(NEO_XP??5A;Z09dbW0:53_A6b\U]+,Z.#.
VIb7[=:F;-Z6]ca6OV&S\:ILMR-^a>V]2O)8?_0W(<=&_.,991B]01#@(9V8\^P)
Y^UQVNTgU2EUfNYJGHLLN_90#LT0SNc>1P;/I?4\SG(<,YHI)AH/F#:Y?aTS;,#D
=:@S3XVN^WI@Y/3\eZKOA898M5?+(5f2C2f:HT0O<VF8CF\.f_[6YLQ>2DU;/gJD
KKLR,/\\EgI<T2a;A1]-35,U>@^AK@e8;BO(,,TcJd).H+#CeSK4AI\&B,0CMK2G
HB@)NfLCLJ>cR84R0Q[.19ObZUIKd^gEI0CF#D1OP<E(##RSI]+TZO\\G0,K[ERe
R:HYB_DZOF0gPO(3P^^.9AMIRd8gB^W&>++)B=H<T:9SKK(5,87I8ZE8-_HX[aGA
U2MO>GS0<gEga2Sd[d#D.U=99]72-WU?=DX3]VQ3.<1)?G5BNM1?KNH:LPQE7D/9
LfW>XMV?KJ<Ifd_TGAfX#NN]L>Sb9:46:>5^-/\/U5A]0MM]=<&?F?fbfUf(cP[A
OAa70SA#YLd(O7PY8^,99@#X=F/AK:Ib?^EMCW&&N:cS==dB7Ha??@7O6V49=?4X
O-:JcfY5_S:>;(K?@ZSa>Q?25C]8TA6e@,<2A\):)V2-/=dgUN..Gc8^XB6YP2&C
QaEbSf(J2HS>bYHR):4d.9<:Nf:G)e8-Q0Q_<ZEQ.EC16VL_CK/b7@VdZ8-Q_AQ[
EFTfQX59.UaFVe,B,<(RT>7O7_Ma66RHd[5Q]D>5HM36PEBEFLGC^A>A@b,Sd;f5
E7+TH3eJ@>L,X]JW(cSW=S2X<Og/UBZ=G:WaH^2-].G^b93-.EMF=R>8J8KFH1P[
6DB,g)HS2/cDIH1cb=C@QT;QX\J<YWCgFA@eK#0W[=O&H=@G.9#[MZ/\CL+N,BAV
).@N;OG/=KgB/748W?EK<:eAA^<UX2LS3;HHI4BI<X6ECYUe2M\UBZ[CeU:KYC):
cB5N]A.D3>DW381R+cWO?&O>+V7ZM40QJ0[IF^=(G+,7:>@:RbAdKPK<LEXHAO/&
b>OQgI8+6Vc;9/0(BJ(-E;3MR\bHWg0.9ZJQAW(0Q;>L5Q30NYgY?C(YbC1N)=]O
DE,\S(9O&\JV.5W=a.R]Y94-,FVSMZc[@7=JQHF9Tg;4&A<bddQN;;,MFB?<FWAZ
;)b4)#.-@&[6VE&b]@B]GRH(O<cO1GQIVfV967&eZQHN7JX=FX;T\NgaW-NX_b7(
8BLZ=0I@_gc=+G@N@PW[fFC+.OYP?949[dXB;.V4_DJ_D,5)GO;6Z386XEeD,:9Y
L5NLJ.V^gM4F0#EB)3fYTVA7JRQAHMGV?AbNJ/TM3VaY3#JPL.c-&1e2_+J]dg@a
[P0=0ILI\9P4Y-+F4[JeXB=<FfI99=Wc-<:.[6dR8[H5>9S:81P1-&@[>]P@D1XF
a<(W>I:,8DV^0@=;ZXC>BafW&(WJR^-(NF,EVUB&PQa<7ATd:EA[Z8ZJ/f;<-W^F
<.HAed&?WS<f,VM>[JN6dWZVDZd<A=8gRP(ENb_F<97KbLY?:]M-88NN.4f=YPGa
LD3:Q)9f3-6PVM.P6+GWI+FJS46H4>JEa2cb^7)0ddN1#I8)OA+EUS1J?@D,NTP6
3[1F0ZVI0;#I?C?K3[aI#?U&+7L^TbI=4^?KE7S)QNS^^>\PM>[W^K6]0GaJV=CC
:>]6(/SWM&0.fNO<S^d4)+V8Ce&_b_6)@UQb;a2d5\VZcIX]CC_JN1T:^@#(NK,C
fE=C0>IC198MbJR>YMS,_S\AEAfRHH(F?==DZAU-D?P<U<VFg,>15O<@_&_D2eV\
-U@&P)=P^7WEJR6+e):0g0IR-W)eSJLKTeXA@[_S\174TGd)=)X5E:_)H<cL749X
<);W,Df47/Z,GV]W(^GGWRc[bPQX814KGA&0]FN(F,5BI)aZMOMWNO,XX2&V4-=^
;e:J[TK)Sc1-_P_JSNO4N,\ZX+40>Ld^X56(&_^&]PF?ONO7@F<^bC,WH[:HaeGe
P_7J3f2G_G;5gVM[Cg((V\U3AO.([+,/aJ#JPH>^^ZVaeI\5b+_Ib?SKd&b/K0A;
4)J\IR/=;KcQD[RUX0(AA@B5\)1RG7V=g)C)Ie]91BH7Z3-_MH<X4\Q27>X[ZP^W
GPI2dM=8.4PX0WgKD[Q]6(F.H54^++R01b_FbMag,BXdeAXY^KCeeM1C3ZC5Q6&_
LHTg3]GZ\;3cB2=3(,,AT=_F<#8[c3+&J^Tbg-\e:A3QZe^BPQUR6cAD..KQZ-)6
@]WIZUJ4F]cF\PPIUL(#0V]15T?=f18Y)]OKbK,>cN[D746HIC.IIM9_OQ?A>DR+
:?MM0E]Qd05NV&I:CQD))W.bH3B[dUHXUVUO/-R?@7U;KN)+R(^KdIQC&J4EGG3+
aKSP:cBG2[Y-a7C<@D^GEJSW>JA++J/3?1@.L>0OIFF>1^AD.3M)bgWP&L4faU1+
8XCAOBK4H?-+g?QO2@bGH1e91)?C;P>]YN=3<CR@2G?[J=H+-);[eHQ]WXSTDdaf
II@IXB7c<d(\;:9<45[4]gC^R^)QOZQ8d/?d>ZXV)95(]-.W>R#Y,)_6#bNece8S
TVL\9(ZWY7#.bU?J9aGB0WUbd67c3\/[KD&.SQcHb,WWJ_&5CR2O6.H1AH&DV??Z
>EV>79g+;PECSfLb]FLcc7-ZPW.\J0,3eRJ,,,ON^?gR_4+8:6,gX[#e.L@O+95U
aFMTFTXM?IRgJ)MKg3IW]7D>(IUAFLSD#aGRW<IE+BE1(dN@M^R)?3VEPIO_K:d_
Of4bV2VHc&Q>9fQZKSa>,6fC59XYD96ZG=Ve+XAUb4<NJI,c+)5NOJCBTd.?<gbg
dR)#?@B^eQfSVJFe\?aNE@>EB2QVJKJ,Lgb,#EbO2&<DFK&(e\PY=SGMRB,1[->6
G;VR]?^(ZON?9N60W\WP07/RZ2[0XO.=\+G_ObQYD2HSI=c88#b&DB4V50ULZ^]3
e-8B9VN?=\SEDFFTD6/T>A53.04+FJI.8KOWI@>DbQ9(f5VYK#YK_,gR)@G6.-Aa
>59/HWF2ZUI_:4f4OS_QfIdM_I7PGT7TF2TFb7WC?=&U+)&)f/E_fPUa4DG7=:H:
PMV^e,MEaF99L3[Q;[DJBagRIB_DLdeUD+9?FKgT1d()M2+aS)&=cY/T-<)^[gOg
(S6#6QW2c>VOc,E1GK;7,1AKdXBE.&=QC[/dSDJ9IT)c,^Z&RdU>MI0@A_Oaf_^e
8GG(R<ePQ,6:X2/:8+Z/:-J0+HdVF5,K<JJF[;a2OBWO6:_O]2]cVcZ],f1VU7,/
M23H\/A,eERXM5eP&Q+>4XNN>:Pc7]MA4.N\<D^&;-0TLKSa4\Z8NWV#\<D1UDGL
bMC?/?FCA81M9<\GRXXd?d<L\[L1^,fSJ&0fG_1T[M:A,[&.U/g[GK\aZE;cF^=X
(/\767/(]-4PV&;__]gL1aL?C+OeQ6)=492K>#U-c[GF>RF_I4JeKg-_g9LO.,#(
J]:bM0.QE,2IJ(&QEY_-8NQ3LU_ac_#D8HT:#=bSY(M_I:T#8KD4:)e)^e13g4H5
0d/.5E@OP7K6V/&^a0(PX]V./0g\4Nc32QETa@^/[K,Z8&L+ZH//AF1_C2#3PPW4
NAeb[effEH[9:2RB^6g(/aHH5D1b(?Y^203/3,K?#?>P_IJUgFOU\K.=RcVT)<OJ
>D=(4IYNZ4FeUbGC4839,d(^<QeP:1P=Z:+2^-FAeZO^#E?;]V[<PI/gTI,^c3Q\
X_dONK]ZeN^3DQ2YZTeIY(/VR?JV\Bb=1?N1&#dF/IUWJ:Q#M0U<Id5d^HBCeU(X
A2(A9#)1Z[:C#,QAHLQZF(6ZS9D\GG5W7_]^V><Z8Z=-Q_g(W/5509eWf(4/]Q@V
B2bD=(IT<eU.URIbO<Rc6.3HE0:VCbcfU5UD>^=B&??Vg7C&U&F<cV,0-GF?J,PB
(;@-GGfOY1b>=]@FFb6XQHN^^4Pc.:a2.4d/>78L?K9SA#V;<MZGa3?Cd5_aOG#[
Y82(-QQgUH3OQG(B<=3ZO_[L]C+0P#[9f6Z@dd#(U^OTE?gY9+7_UG3U6S51&Y7;
U&d_:JW[T25H;=ZOfP6WZ7DgOPZZ)bdDWNTA8(5LGbUG;#8=V-&[DfV2NbMQE<^c
aU<#]J3,L3WYB>@C.K0G2@eB+;gfLf1S8fddfR0PWXcUKN5]a<)\HEVK(9WbH]H<
G5<Q7ce4L7LJ2dTML--<=Na&=2CZ,?U588JM,9;?T?e@#ZT;85HXf;gQ97EK,aS8
fa0+)KM1M<,Ngd4JaZ6[NNQV>B-1J5(d0KdfDP)aKL^G<=#Y4X1<)5W^<bWOG8-+
4,cAV+a.MC[O+b7,SZ1H0?b#+MECCdR==W<af04V7Kd:_14E0f@d\:)8I3S9?)g^
D.J&SB\D;Z@QT[Fagf0,T?MKPMEDWf[?/2\D2-Z^Z;)V/W)J6Q#4]cd9[U31WO)c
Z,B-f8VIg3G8Ag1@^<9c2?MWI+HLS7<faYHUd>gHLcA58EX#HcF>8B>Y&[TGc5.1
E4X/=,=&8?-XQ2,XePZV.7KHUL<aWb.#NP?g]?(?T4+(KNQNf^gSB0&^7.>G17a/
_De@@fZ/C9_KU+3-KFIT6Ob/+LK4TF4<Wdd9VA9;[6ZXa\]6=.YC\?\YWVdgZ7-K
Te_[cW(@E2YO@6:A4?&]57c?/[A3KB#^QMBdaM<0521c1F--a_A\(0]-)]CJ?VXI
<&Z]Qb;#Y;[4>&6I#W/U3_,33FG:1M5<T\7C4S4ZI4A5IP9@0d_@ea8<6B7UK+=E
PNZYO@K8&]AVcI.1;aPXP;VQ.-SCOZL2,0F..6Z;GCK<Dd>C2I@d[6a[)fV6d/^Q
;;04e>OT@3UO@.BZ+.HXD>BGK-6H8)4-1X_B6R\fG4c:Ne2QbS]TgQDE=I_/.G=8
52fVPQ_b,:Q)OA1L)7XEZ]1OP/bOLb2VDVDKeT@>39a^RCG(O\M\@FgeO2GRV&-?
F+<V^[2@-.>_d:Xf,R,Q^INaLWb0\@cc(NW(F;=3ed&Y:3G<c1R+HDUHK&:.a/Fc
F<XdG0C6ed9@a)\5M300a+4[dGLTg)O8+/IPfaI9&64]?2gVFX:&d/Lc\,1[153c
KYM0=45]@<.^>M&[Y2[;4b[IB=?HBGLGXCeN3R0VI(a#a<JMN8K?.[6?0g\#@/#g
38;MGJd=U^<W_LIBgDOD1I_@2Z_[/^G^;;N^87(M1>EgLgH5>ef#9VNB:;c\?cgW
\:PQ@Se#G;=](IGX@#c)Y30/aWb\a-.QVAXgf6:SI7D5;M(P]D</@KdUX>?.]PW[
J.VYL6OBM.0;9eYNLJ#WGG,f@<P_:NC7UM#HE+-+QeCII?6:)O#g)R;KJJR=aJQ)
KF)Q&6P2Fef@_[^^X-XI\4Cd7B7MdI1EZ?HaZd@T30ZD1U(d]Y?A7e]YfLbW[(S&
<H[K0ORCLfIM)=K(YND.]645f4DDV@SVHa^b/^[Y6<-N^eUD:gI:S&#F?aP=]#K2
I7>:\6E^Ge]FZBd;4H5_M4TK3Y1NQ9+BQ?.>)R7/P;2<3\GOU6g+6_BTR:^Y1>.T
)#VU)&ZReFd9bI?-2Q/UT8KgQ72_WY3E3Y15NW-T56^4Ab8\.e[+@@16g_b8;E\A
][GCJJP?aYZc2I+6J_LYOdS4Ha;HR:)<KEM(GC;A]SO#U)a^M(\(T[G2R++5a6>#
a=ZUe_KV<-XK?1/GI1?-Dd=^>F(b2Q8R2E>H.-<1af)HRQTLP:T_fQI2e.EfCF[M
75[<?#c)&,Qa^\f:6K4@A(R@WXP;TAL>)a=X<f;3)Bg@aZbfO397HQ/\SFcS&48A
:E16^YXHC3bf5aG^G=OZ3@/:Bc>K:@-d/Bg4/g+2QTfY9/;O^.,NNb_2Lf\3+K#<
<A?e3c.NU5X;3;W&09a0;H3O1FadVFS<ZDFg7IK]WXCTW-IJIAaBf22a+6]V^6+e
@:GWUJ-M/=UQDf[22,\\8b4[>)MNSDA?7aYP=a<[[(_9eg9AP/bG4\S9IFJNZ=@<
,>4O2QP=VK6F?\^&T<S]N\HebK5^.45BY+VS8cLST78HKCHYVR@K_B.2eTB\@bG<
,\Y^9c@))S,Y&4#fZaS/FTe5(5CW/TBFB0]?b>Y/_N+(H);,J&f\,?FZ&YPH?D2\
R?eRc)a^;<Q,=a&_0fPL=DI7F+H3X,Q5]V>gE)A-X/@:b/>eEKE]KK8Z9UOFdZXY
R;JBMO)C^aR0P@,0Y<Of#C/6(&6?aSgD(c9eB7I7M^K.:QKRP6+C&\\S#6-<401C
f9-L>:KffAY(d,1^@La;f<TP[EWgDUSN<.UHQ48TUH5DBM,F=1f\18&^<RcbMK).
+/d9+E?_gIaN8EES3)J>X;?#I=_+VOdUNIC)^]_K/@YIX-_Cf>ZW[5D7F:4)PX4T
C\X@5E4=<-(+@Y(U2_)f16LDd<eUGJaETFT;(H#(W3gDdK28YESb9NJPX>#),&e1
@0S5#QS1-FP6#N=MIA]^A=JX@B2UK.e+P8d.[,S65M[:XNI\;a=;?7<D<H+,[HOB
6gGRfV=L1b8ZR57NFCC\7G\4HIfdGG(FP;^XQ[N?83A[:e9J0NS8YaBK<a8#DXV^
Y,OC>H^CX)EUe>&eRg5JW=X-JfE<;B6B,a8d79_eO>.6BAFL-_NO4<O70FD,_Z4T
+ED14#+PS#.bG<DO[U:g8#b;2bKaLb;F_g_F=@@O#1f__7Z)SA1UgV+IZWdBYWGb
Qa]DFF>WdUg2J]KNY0DR6L83b4MTG/TA-&^Y]0B5>,2]Bg3E&+=+GL,f(^I@RYM]
X9<8cC5^^)YWSET2&:VUEWLXD1G^FDO]g\(V19O[.CXg3T8e:IUJJ=IVf\Tc/8;9
[PN8C38[VfX?HaAW7AD:4?Z)_/_Uf-T_(/0dBIWcX0RN1Q]W;aBENb1a\&:6R#CQ
-DCWJS4E.&D0N[bA/OSG<5DA5(gL:4JY>NAA>g/D5d8fZU_QRJ.Z]&Y=a;<T]RD+
4N@&_6aB&cH2<=EU0EUH(EYGZUZ>QG2+&E5>Z_OJ\2g;13SJ]3JB]096a]Af)^F[
C@5DFXZ7Bf]V0]JU[+XJ].R64=QLD#Z^N&<ZA7eF;A1eZA\<:PNO)_>B#UK.W78M
&7(@?\+&eK84ac2gQCIUZO=DJU]0/J:]WVffI]3-:X>LJaCgM8YB]>,M(L?HWN10
.H3=D4\(K<C:YOe.TTXRBDON\#</)\@=]C@d.<N?L.19#E,+G?ZI.__V9a)#JR?8
B(aAd@A4_7^[0)Z=a&B5+;H6@bQP4O349_L(,6WVKc8g:?UfW?[5-_d7/6:CJV0V
?SZ6b#N2ASSCX4UH./F=-V>YO\@g,+UXB-PF[3@?78ED]A64-Z?e.4_OAE&4WN+=
B06MbJ,SE:b<\ag5Cb^&7Z]Y/U&[JMfS4API;[aG6LGR2I?6Z=_Da@^=b@#?dH8Q
d4RXYYKgGI6PA2fEAQ6W+M-B<AA:cVG1O@d=6SScbD9,fa\HJ_P3-[V=TU,4;\Xf
2VcOG#8,(f.F+cI&:-FT1QV,S(#<7&eTgN9JQK?LLA;W,_#U_G-):E@A\H=ER0L9
@EUKO9OX@eNWXFCF,9I75g^daGW3@^eg?O.bFM=:3#)FULA#GH67-B;J.)8&#ZI7
8/ADT+DO9F6H3(997+1H^G?3<S(;QD.R1SZ3X2;9U3DL8gDH^(N]^Q08/C8c@g)0
D)(6/2_gF?SJDO9ED@)5?:^H]9=A]^JcQ3)9YGa;-[=)P\8=O()M-(D[3eWL?Y51
F3-A2XU0WGW6e6A&KMf9/Z[];d)9NN]O&b^.2QT;c9Wg&g=cIT+R#XZAf>Ic0f_O
10E04UM<.I;_^K=C]N3:,I]MQ8+>U+b6H,@I-0\BWXI2?,+6f3U-AHYO,/,C\5.A
5O51[\d(JO\VFCV>NH1Ye\FB0QP^&7_C#dC)fJ+ff:gUI/J\X\_KSec/^2g5QQaU
2d/<?.UWa4&<T:Eg&g?3UYeXJ=F=R34>\<(63BXTGH\Q&17]3776fS?7;3&1GZOS
Wce?fJFI>&]Y_BV7?./ZW@^c@g1Yebb,(D@8]gZ<L[IfB))E+Hd]K/CYL,8JO>8M
aZJLe=?Y.CJLIJ9GY8WG0S#3CU874E/P_>ZKN(U7;=^E:W.<Nc2dgaM_EBT2A.,E
/:ORE\T7Ed_/c6<XDN?_KSS?+9e@:#6202OA86RLK3<EbZSNe53eXX7P.Z>,8T=Y
c1+(<f8K-b[WC,33VQ2=6_8=O4=aUPH0@(,Sga1]9^E+ZaUaRF3MW3#<TXU&42ZV
9F.3HC6bX9ZTCI#a1[H#e[V^3eJOaA(X;R>1<fWaO;4@EA>]af+\0YU54<gB1)7V
\IDGY<Q9e5]Af93W>QY+A1f9CGLG.=&UE-g+1,0B.6P57:+E^B/aEL\YPD^KECM;
2L9]1@D\c\VT?4ZJ5fASf3be?HQ]UKKSJIfCB/fPR+HPB^Z.?R=7PNI1V;N>PSMB
(Z:ZE<QE8UB(eO-N\FM>H]R9gUEUa;FTbC<WI;BR+[d7c+I8gSB-P#:g++LZQ&(2
Ie+bJ;J#WA9)XM67?97^.GO5;<Qe>AQgFR[6OM4f)^J]AZd1GKA9C6+V^GF)d)A5
gCV72gKE7=.HcGdgM.R+9CGG8861Va6-HU@LHVO=#).\N@0VYeEBR=0efOF>,1P4
^U,Z&T\3A.6=:OW4;D3WBI7K.OT<JQd.F17S:cI#7N)5QG^_6HXFgI^P:=M-b8,-
T+IA\>fe:461D8&D>E;-]+_MO?ML^5:4F&[+V:g.6b/)=A3L^^4?6UcDJ>f#:B[<
ag?;bD=;FB<3-3c]H[PUEHbRLL5P:VMLO&ZeW(9)bff2^=[7,B7HP4P4ed/a[]@Y
0-^8[^976L2[/>R)GeX]]XF^6+U<bfY>)Pa(f_fZZD-Xa8,=(GJ#\=g,2<Q]#E\P
/QGXM7@5>DVJLF.9e68Jd:SA;?4O>9^T4)Y9AYMKf&7C<A).=;#WRgO.3@&&_P@-
HE5:OeYQEXCPB2,8]GK&[WISa:SU2+@PNQYC\aYVQHH\SH\13(gGNd-)T-<^6g/E
U_M2f+G-,T,3IFOMe]#)DNSOJ+N)T#7(;)+2VN&04Z?c+U\.=T:JJ<.NHR-^af;6
4RN=M9#d&FNgJWg,bUN7WOCfZgYX:;X/BYT4b]8g9+U)N</W,OfYZWeGJ]KGf]7L
H?S3T3#O7\9OGZ#K34#f9SULQ^bd.e,QY=MaIHAFZFCZfUWH4GR9Q6Na3UZP]a+S
c?b9S<[^ge^JS5P:RTW_IG_PD?4:XL=RK=fG651SB?U;OH6(O+HDVTF^-DRN[+I3
XLN?>3e_VS8,(WWC,EPd?3_0Y#cWZQE+dWcOWT.W1-gcO[1?T@J2G]gIFY.EfK=+
O6&A^T8b<NY7&bNWAJBOX;\+QCP9N15&V=7Sb]0P.]&_(5)3GJNG)Md^S>fa:UO/
Ve?.<?]IFKZ^53b(7M5GYLWU3BcYJ+B]X)5SAfOHT:eL#1fUAb?I=1=CP)@d;Hce
<FR\ZWVdH7F5=^+)P1[ea6DFK0+cV3.+SI@I#X\;-5HGP/c[AO2c+Q80geC=]1C=
1Ca+4O#6.<H+R)].)/CLFCTIYNL8Z.T[EEWK=LA]2&dET.5S?7J:\Q6NaM68E(FM
X<S@cI2T><?4KD45QNRD-fS-TGPYW6X64g>]]C@5a<TVFI6-3H,XLE5WV@?#+KD0
7.0LYJgHIE581J1FV4LX]&VM<=WCbgCY/9b8/.dda<J_,,bSF6f-]MQP\aE2YUEJ
=/F#)+aGEHZ4@B=Eg.7_Q]I=5]-V\-T6GC^=bHb5]8W<ER-S\HJN=O#cT)8NSE4K
[UQCg=:^LS=<DB[3&,,6I=8O+/P-QJ6YD6Db^b.@M1J(DI^^9HIN787b<Q30.1eY
Me^LCH#:&;?-9)5X#N.]caJ\VR?f7CS7\#3B7WJd\CP[2[VQ,@f?\)K>3@#P_?/R
-/7\TO;T+1XF4d1b[g)3DDSUd;W@\IK.S37Q5:F4NHNAS,<]gEA90Y4Cf1W2+S_3
ZD1=JKBZSe(4],-G>/1RESB&fN3#DD>OS#E(,\3X),5Y3YH-3PE4X(F,]I2RZAe@
?#Rg-[<MG;,(OP>\eFC_cRGWX>bKN/I8B.X(CIQA0NZUg+bHO)28PUM-VcZ?eR#4
U=_XDKI\c@DX@9(2GeNAf9AK#L3<?Q5H[/V+G0OAB]H^6I3W,LQOS3ZG^SdSU[cV
(cF<EX7ZXR^-DR2D[We=2cM-^-M&.SFOKGJV+]BUVPa\#d/#W,gLSW&JO&@SBUa8
:4<G4,Q843@&-GGF)^HATCbQA20=Q;9TfC)-=-Q@I6d;?7GH&L[b_LU,a4LL<Q5M
FKa\M2A5HgW0I\:H:L:+4S4^?e1FXTb_<ZJ)E&TJJELAKCf6;L:,M^_5d<&KZ_TD
WC,#9)0RX-WPTZ)VEQ8VdP7cAQ12ZA[d,PSF#00eQQOK_-d62QV1\AELR&>D6B+6
VRF,LY+P@;U(4M^:gZ1&JC<KO]<>2X[+045)T8DM9MZ?]e_R7-&J:DF5R8RPBb,:
.@3\TNW8P-Kc>F&L8UZ[6-=:EYL#:3VEWE?Y)1@N(/?B\=)+(cE@YS0)=5ADAg)B
D&>-NW@P:?>(>V>.J1#Q^>FC4A[EL=^AJB92eCB(B<G92ffNIeUcbZdUU8b.-Z?M
ZQ3IW5>:K\4ZP(>FB2YYg?Q=+,AZ>-=G3Pa;F-de9MbM1+B&Gd@5UWL-\(g07f\>
DGU]LcG,N?dEX7cYVP(NK;ZK^J^Y)>@ABa?;P,E?HA9NfF;\RU;:B2A3C0^<KKZ]
d9e3:d(c+]6+a_K4T5.Lg)/T9--@b4?#9fD>&DNaWQZ7efO(63Ue-G,^NXaR4a]d
VeRVLg3ff9-+=I5VI_5VF6U:.cMOV=ZNM>BIT.,XJ0[N/A5OSCeN<\T<I#VJ))]:
:C5LO)PIR7,B#;Mb72;/HP&-XCWS-;><SSf^</)HP;4C1d9;6I)&KB3&^>?NC8Re
HYRAFDbA(/1a,HDAD73G\Ha..W7J5&e_87.IU#J4#_<bDWdTW5a^X1ES#;4,gIR\
_0,-,,2,I^,^O\14?9dRMW6032LBX<6b#/3B2M;F7O^//Z)156RZG4_D.X2L?KOe
g(3>?#((.0_P]eb0O20@&M;SbUR,HGgA\eDTS]9:cg]R.PSY30:HJQJK?7K^9S\@
RP/7aP^,NWCO9c?JS0_D;ZFeSSDEb=g?-QcLASb(ZcVKX^8&cA[QF2ISQ#C(/f^8
4N37S9Q(a/\7F>9Ba)F8ZQCVYIW36Wb=YXdfKW+Td6U,A#\0.\,-6)3.g7L<G.X8
V6XEBPX+f54C1/PdJ[.D)T+&NJ(R57E=eGZC_<U385]=EbFA47L1&/DF2)#&/HMG
&W:[?S(?bW[Q\R.,APgMe;ISM1_82Td0U&S,S-^8e1PYNAS.X+e.Bf4)G]d:<8Zg
.;O)WGKB:(aI=MI4.CL>G6L28AgF-208HY2\4Q1-D)2K@ED=d1.UM@P[JYHI(gT\
Fc+R=BB&Ld]JD=/F;Q)8/)?d0(5TY7-<D)HSeVgDZ.4K93:J12P&+Y#UWfQEB::=
]39,.0=Vb=Ob9A9ga4Gfd1.S+K3+\\M?gB7(NeB#^HgL\X/]I:c_0=@gK+YW?F]G
-JQLe4U07=]CBJTN&I\,4aTV,X&N@PF^GD<Y[REQLfX>e;H@GQB;:6H-ad4WYW33
ffOPQ=5G\\<W,A&JRW/g;bT\YcfF@/#3F:=W@+E)9O0UcG19dZ&36U=1<,DPJ]a7
QQ(H2@1K4@SQJZ-I-9e;HFI;=M1PY^\N4M->LADK>5-SFWIW3:_#X\c0Q,T(_>G&
&CO8.9PM@>3F.:Q:_N#\GJH.+8YV.+AdYaXB=O/@#)1Jd;^PBJD#\aSUO+]1aH-a
O5]^0HgR<Qc1=_QG/=2[/,P#ILUeWVHMbH#[b,I[W=4f_:H:@37RXPUaZ9M_g[aa
]DQF(,W.4KTZ3cZ3;CR_K,QYDUa5b&#7,5B&IAS1\=ZVLf]Vf==/=<6+B<a]45>U
VT^9[QIU@:6e.1+U>L6Y<aA?BL[DG[7LEW(.S2a2XX9:)4=VC4,d<:_-;X:&]5fG
5HZ>&_d?Z^VR:ELbM-e1+^aO@L&-XfI]L_Q5XcX^T]E:_;Eab<3E#)eRI)<bJ<SF
<A^4NT04FN-Te#-@WZ<VR5ZHD?G..HSIP5<>5=#W?fccCQ4ZBYb^^&RNL2_F([Xd
7BDdO-(2+KB,V,DKO,29TfU&AR(-KaN;([d(\=cI/a,1FRfEV;X8XZ]FdYA).KP0
PQ@feTd4GeC4Z&=Tc.cbRNH_5e>;:7:=O/6D3#fU\9I;#BV4K51<GO&HUdJE3:dg
K5WEWV5ePS[M;,NZ@M&KZTJ.7gGF<M?O;9,C,KXTZX.@9[fH][cP4+<V5#PIVC//
Fa24VY7B>=^#18LRU\e+<F0REBB#2E\OY9dOc?0Ta]P;W\8d?7:3#8gBTK\#10>&
d;YO66YW<>@A;Q:dN=c>^#ZfLW1]^3/N-YZ9DHII880U_8F_gJC?b5^1(-#]:>[A
Y+4F<V]#+A#X[DH0gPKb[gQcAZ#W+LgaA_25fJ2bEH4_:X,PPEL8W2QQ[&+\&g1J
^WAXU3Bd827.KI/f5JK3[_bX/\\]:^GfW?W,,2aR3O9RF[/27G.RM4NJ?bBg+WX6
>.8V:>d;1/#HggKTE_ED&T/9?SE<[@E)\aT[Q7BcB0J0b279g];e]R5;+UI@8616
U[DP1Tb(UST\83_VeeRVQ:0EZ4J(gIacKcYXaC0d[J&)=#TBR#6.Y;Q&Z.P[\8);
<QNWOFJ?567@G_AU4c,8NS2G_?gI(_>0EF,I733Y;XJ#b]gRHI2)U0\&8Q,0>gU1
1Qe<cM5:f)U;;b7Tb:N&:=9a<)-WT4dcO2\X-.XaP)PNX7X2KQf(fABI4bHMe^_Z
R^Z;/^WJd:bN&^RYKUZ\/bA\M+6ZbOPQBF_Ef>SeNDSM+;@.OH_6JFKGA-[<;-A7
SaQ8a+,e,Z<[RJ\KRC+\ZNf8SBLcaQUP5:-LM/B;fZg_X:B&74WBGfN(OF+bB,>V
fF_II^bC6&ae8e\PIV9751SdTE1QWP&MU&OZ<K+aG@YC0D-b?\B61LE,;UMb4PTX
3^;=CORf#QgV/8T[/XA9X1KS-D>.VJR.g=+T^SE2;@@]=2&B^6//3Y2B0eODH3fO
3/CcBM^0gH^Fc(=4PW&bN)YKW6&VcHfW^\6?S8<.>08NY0b2?S=D5HJedSPGC6U;
7>^BZc0S<gCOWI?KCF?>P7054HaSe/7S70-EAcB(eMWK@8c&OZ<<eENcC#Gb3^.\
fI/e9e#ZJ;&>H^3E2>1bNe#5Of>+F(9_HWMc3?=[.>0c^?^.(9c3V/HDEV[]]8?R
[[d,>7N>P.]E54V[eBD]IV+HTU^bDKfD8?-RBY<Z-,73OdOe-)gMdIK:0K<SO/6Y
A/,NbbAdE_ZK@TJFUg5NK46LWHBbAc@C]3R<NH)@ff\-fGe?b=R(A[+Db@_LbfgB
:OOJ,ba-f3/+R?D=?J/+[+GM+&59D\/@LGPQ,NLP7P/>60<=_f)CZ7Y_DXP]T\UC
<QY+\/Z@,(8N-U741H,AGTAa8,[LINg?Ac?/VID#5MKL2_E6?+U<I0=@I72]EQK(
><5bGVeHCI(.51E5=NVbg0H/-7P6=fB0(JeUI)f/_4f0RdcCgVO=T/;MAO]667.Z
IbB^;602W##fRX-e>CA&+.G>:Y&NY;cN-?g8+\VG,R#JN/50);Fc6NR39SE\)e&K
]:AG]fD^CQ/?=?3R+<#?VX,Y/OIFP\b8SIHYBU@Ng;-6/31Z21NfZ1V#O\]cg?f1
UdH1K(\?-d,2=Z5-QXaH\DFPd\HNE+;MX6JDc/O,MF-CB#>G73X&_XC+Id+fdESV
5XUd77K-SP..[.IT[2?E]VPNfM?A26OKGX9-N#e&EEP>e:7G2>/(X2LFb42V&JgK
<0ScGV2(;[FLM#;eVe<.-IK3(GW^e&<X4S8B[?N&CXP5e8@89;g)U2[QdP,TA.7?
?]X_bS08F=A]2?^SAYN=_fBK=Q8,Q14(LVS2-E+[C<1&Y)Gc2@D;?RG>(SNPZ3F+
fWAOC)U>2fg,=\WL-8BZ_X3FY257,F84e]bIZS=>BP\Bg4=YBeLMg&O30#2-OFM4
gfX&?[Y@F6V^LfD33P)//>=1>#8/g?_ePb\.U#Zc+fCP5F2FLa(JgIW?M>6VTR?4
0e03SbgaU0G=B<@-;NCSDXX.Ka2F9BYPC1EQ&93aYC[XZ4E:C.V,GTG8(.L&EJC(
2B5,5BM>;-c3:L(HFXB<7^UNN\L#5f7Q#&P)8]86NBL:54YVK2&5W4fC.,G1VHJV
0,6_#:R5dMH]:LG-J.(Cd-8416d4BA5/?09]5^<[FS\TO2L\)Gc.8IL.H]B1I#YN
@+g;Z)d9?@,43e=NQB:AXW\/;@ZD09CF6#&L>7[3c?eQXeY7I9HYc>X;cAUNBaL9
(QS9__TP(1LWZ7aS^310aQ2Fg[Z3bJ(Q:D9,D;AI/CI/3Cg)<>0=DNT(K.5.]^SL
;+JHTa13Hd?F&V>[2dBb#ME5NHd?-G:dB@f.gV->K,8DEe9J,CQ8Z44)ONG#;C[I
QNeR,K]=2_[b2R57A3^)V.VfN#U^QUf1[2(;;WE^efW2#A7:)O&S,O3WXTd5&ABN
8NQWH6)dZg8Mb8)R&YcQPOP:5[-:MD1+>SeFXgJJ:<aR<VWW0a7S<PVNb3KcSG)D
Rc.;0CH^0f)+:T_ga.?FG&@EZ-:V_RW9&F77Z0#69G/CfGgdRFE@X,6QKLBT,H?:
g(@gfgUU@6c=e(LUBV&^OBY6].,EW/;]94Oc7=PdWfeYDbE3/dgUN9fY-7Y/NE#I
V>ggRDO2)D_N\30cPB@O102)+@VF570I2d95(E1bd]X];V=LJ[bD1VYN&KY2R&R5
OV/gDS.fLc,SYK^#L_X;I-N96)H_?O(WS:U2D3K&_E>fb>7O4MeCI,ec0WcM)2cH
c84;J#M[BP\d=cXZ]AHDR05F-V[S->2E-U/L+g2+XNPNY_B;#b[e2FMR2&H7-^c^
3D5@6A,-&=(:Q?Hd90_/;DNR)JbETB^)XL<VV)Xf0/-eWD_&NF,0T00STDL0)AF1
7]X(d#PcS/-Y+Wb]\A?V8\JQf#65U8gG8d=3+g)>IdTW=TBdAIeU@UdNG^TP?#a/
MVeGFaX2?[]]Rb\GDT&AYHRe#&b#I:,c<@C?[,LLaQKXQ9)J?77K>DHY&fYMBOTR
Y@F[W/QV)cFQeB5;e]-?<B<(B0g,[\)d<BKA,^D;\BEWL5YR()S;/DgdW@W3ZMT]
P58H,aP3SMCa?gA?83L6c^\7T\@V&_HR,ePcXG,L3&MF[4R&X#_6>bb4_1:-f]GS
NSFUT@00IQ<TUJ;aANb[@^#<;)@]A=NCZB1[cP5C;K2U&e[>=_2RGa\\]fI(T&HK
#@7G\edd5a?b[/+0gZ;QG_RQ-<)3PgaG?_-f-@K>LB?&4Ge\O^&2PF>dF\6(P6?O
&eg,])^.&;X_L3Q^G7#S;9RR6<+G8+gOZ32ZA5/Ed91NV70,TS\\WH=fXF91_7@_
7ZE3^_YZRVW[UNYJQT:(^U/SD)ABe]O.X2HcQ,\M246@8Be7gE^_=e[-=+YCPadM
@e?JD>)NIZ/HO4]eYMRU68dTU(6FTT5]@)K;d0N;IF?P1LbU6KN9(c6BA_4<Tfa/
.8f.W2MS-f7U2R#L0/=fYdCB.?ddHNX:?g@U21=9)74PEZ7B@/91QAeP>T?NLaJ6
V^GR\&a@KV\:LM012Y4SX9D=:&ANAM#8F?79X&\Gb+;9B^ZI;5e]#,RSa:T14^@g
gLRX?80^X=_CS)b^A/?>DCA)=E^0CX=B)ZBb;_ddLS39H8Q^b2^+Q4aH_&I2,.YW
Y<=PTbaYN3.KY\RBRF1S2LE]CIEMV5EP//3Y;0cW.OUQ-8KB3:S&K4]LR.;IM(^7
>QU6\?V-P(+B5.dS;28bF-DLJWW7gFB;K)K:,_C^EA+IALNIW4adC6T7b:H1MJ/W
S&_8A3cX-,./=4Q-\/#/0\>9Kc/7+M5D(&&I#,[42(-/O<0;B3A4)YU5g7RCT6TY
-)?>&5H/5S+>gU6P<(,Gg8#;2C]7D&3SKg67#(cbV@e@\[PIE&@&II<E5LCZ4I-Q
O<cNXEUL_A?TC2?>F3==5S\\A;P^EY#9VNZK:fH5_&8?W^8@HQg?_6cFP-6cScQ5
#A@-cF+]1R6DWZ94]a^b76;5b:OLH:@[]=2Td<02EN@C<?CO^EVR6Qc-:>0Z,#gW
c)WGVQ[7R3#-(TT4Wa49@KC;FZIA,WU>b1-R^Mc(g88].FUSPG&71C=J[#X^@T#-
NR?E7^-YXgZC&0-G+]]RD76+QKNdZ2@H.U_Nf3D-H^QVA8D#8A;](^7B>_[WE3GC
IB=XXU9<\A3?&)^Y74T:GdHb[B&T-RRI<99Z/-\RGEc41.<KYMCLSLOe5\6;-f.,
O)KE7&^:(,cE?]QVZ+J4:LX#1^XX9K]G8A^4C:IW+dAQB0Se<CEQMXHUT8KOE[^Z
Gb-[gB(D1[T;B]dINXOE?gb>:N-?ACCJNMTS;X7\gP8=e#D>GG(UdR<:7^1Ccc76
#(ZRTARLN@3]Yd,SdRII3AgG;>?JgFM\8.52Z&Y=FZDNCPKWFSce:?@)gELJV:_8
4HZ)D;:,7F>YYL(\:&.6S[OR&(Z5PH^eP/2A\5TCASVNe.E.6?(P9:TAC,c8d@&1
7/NZ;fGEV_V_[)&J[@B(GM&R<.1fe3WR#cO8/5:GG&4eLFJI-YHQ555+-W@ZI7;?
QLZ;+)\57.9?@<Tb:O<VNHSVa06WD;B@ZPM8aFY5.#,6)-M;JA8aVB5VD@@62#Sb
?a2+M/QR0dd8?K9JQ5DDdA>>WG/#&[-;PCGURTZJ2D-S1?E@P2/]2:c;[D@8d:QZ
(e@Lb\_BDQ#=8(eS0O9E1KV]DRE,0c<<@<R+&GIaVHKG+4Z)V^a<cU<KKb1W-+Pa
:DCZ58XI1M;K]+UT<34)MT,VE7eB?&[?JPIX2#fgQF448f4AagK>.]O^/+AMC.:<
_c,T801:Nb7?c[.,+TJ=8JM3F8FUHeX6J\QJ[RdP-BB\c7DP9PRX,I;,8RC8#C=O
4<SPYU7MBV]HC]g78H#_44P,&MR^^Ld#.,P3&::Y3JFGaRYf83M4V]Yc=>Q,U3aa
_M=MEO4K62BP-&=C^YSNTcY4QS[18(3FU#)\<eS&:9HU6D]dXV=T[;:HdQ9?F4:[
QPD0CZCgGOU-V>?UaURK2A)F2G1(3R^?TK]R:J5/C/^Kcd)ZKV-KU_^\[X[D?/VS
8DS)=/N^LA4,?6QB/50S]=C+a+T;V9Ae/CdcSW>LGLdG0cQV,4690/YI6d_aZgc)
6Mc4N#U+_#M)HA6YG,+&?K_LGb5gJ8e&+ec;Y-/O^dd=^<I^DGDX>VG58+4(.BF-
N1EfQV#Q;[E>5U-UJ+KZU[)GDecUJ.cPMH8D0-I7e?VegXO&f<BJ[.VW22UDb(V3
GD\.OV_-Oe9RUPHBRTFf),?1M@W[^ZUe3OV)c=]EH9bW/;cWdNGHPPP#[VG/ESJe
cN6+bH)5A?U&6B?G4UfFW7M33<ZRdK[0^8gdeY5.4492ESD\c]g/?-/UV)W3Ga=R
SMaT&360#^g:]LJG4d)4?B)_5Z)5B4BMg6O,3(T#6S>PfYbU)GNC-4U2<6ZR#6DA
g4L_gW_QcG-;PH9I_+YF1)(HS_SFed@3VOXPIZ=C9)^TJX^BT=#^&12>@bU.6]cb
Ba;d3Saa?5GJ6T&cWQ4KA.J_[;4<&G-1c==S9&?S8E4d>5TJIG.aF=^GN_6MUc)3
OZAQd7Hg6[RP#T-:+IMP^4H:O9fa#2^Dc;.MH;D7XgR6Vc<-8aKcgaAJR/[/-ZI/
dXU\Sb5d5-TbGG?+0+2f.^=IKV<=GK^@X;1;RbR&L-GCH6.R@&CP(H,HJ\M4?=^#
7?aC:e+P-9F4dM/M^GdO2ccOM@SUcR\M8X\B+DA<BA&4B>+eT3Ua_g?AZeM70gR_
F4bD+A>f?BN,Q2cM,(MDbQS)_7X1/1R#V,E.WY0]+IOaL^/<S]e05V<?E,LPVLMS
?@UAeB,b]HY++GE@0>cZJ<^eReAW_bP8c;I3-BBdA]VaV&9RC)-^?#;N,SX6Z<.e
RRId/UaY1TE1fK+Z?T7<ULaSf\V@FQYD]PZ/+18Pa-fRaQ/c,-aDgL5YHEB8[(),
>bCfDFEXP.NF@2JB(BHbBRW6O#/aa5H6QCUE9d]NcE2QTFUaa(^HfKg1OC.g[XT1
PbFJMOV\I&>3YB,RMe.A[:^2BXd.E-dfDd5a+cR>Yd)(<?CZH>b.]07LW>)99>?H
AL6U4.CDWL).&gNdebd3:JS9,9UN(X)PJ4G-[1Mg+YV)K_H@1c-gVa/6[VE7I?-O
4fb;.aE9KU4(KG5[\VUYA\YNRFHf_T/RE,Z5M-MY?f0ONX6=.J\gQRD<;4S8d>M\
6cZLTB]0GYT9D_TgcF4aGd6#M-Y+)X?B<,JPH&[H3P^MJWC=<57a^>ZFY@<d7Q@Q
MdePSY?UZ?B2;&A)QL-M=gS7fA-^d/_7RNPZ_^.JS8HBXb(6.JV+V,8KHBJGFKKS
&9+D;B;Se[XYK&@P,#QA/LVSCTbND)cLM(XZJ05L<SQ:)b4BC)U9.3.6FF;Fgbfa
Y5IbC))0RC?EZ1aYRVgG32\&Q[UScA&c-BO_0T@-;.L]Jd(/65)IWW3]@\@9;@<a
B=XONO5FCHRSeX0Y6.e(E3H(.Z0GB84Gd>A\G<\9aLO)T05#PE@,F;Y.=TJ-X#(^
ZP.;_bb,Kf<[Z1R^Z3)K4(f_\KB/SNNQ/fg@?GDQ6^5Ka,d#2;7E:E^A^U;&2\a@
/#Na[YY+4+9;7edgX6H5[R<::-C4>QUM[0]55,5ZUO<eP4f]9USIZO#(O&FEf#NU
(@b,+/>I(XF@8I#Y-cA+8V:Wa[):<,30,E<;O];B#0KK-c_WN1<#74:JdY)d=]+a
9;f4f89K,A>YPKXO1&YfVYRfd6b/LVH2W5SNQ?U6ZFIa2]K2VfL=<<\^ge7KE5Wg
dSF_=&NgZ@1<d,T[[+8f\(@:c-;)D_&3#ebH(K(9g)1)\-6//fg1&Z,2^X2F5Xag
9GADK/b]Ba/B?#6dbg+?(M8.D[a7H:FKPFETR@[;Q#-/.P\+/EG.He/#bIX>O)(d
]R0PPX9HN-e=B75#Z-&F^d0c0eML;T[PU<:,+KQQXcM@=SU-2ZDUF/@ULKPWC39d
a(Af(DLJaHCFR\\6EZ1G;9Ig1LJFF_K2O5H72_(20JbM8PAMH8III)S<APTJHE0.
[6C<&ESVZDJ4<2N;BC:@^-)Z5]E^V2.,EEAO&&#I(?F\AR-FRAU3fVcYIf6-4aa]
,YI^HG\27,d3SC?Zd,&P+7+2/QT(>H0ROQOTI#_=/O?CHG_PXaU8a6)1<9aE(NgV
T<0,C&9ED&H+H4.2]@_aP,.GJa=[K?UHfCH)ZJ,V(#>:DG@A\7(8@c8^()BR>UE0
5FOgd<U-[[9HS7QB7>^,CGJ)XZNGL&D8cYM/<\d?@)X]5UWWZ9P@3)O0T)SfVUAJ
T+MD9ODf71KM??Le^PUWQYBY3&A0XPOT05H[TbLS59O6W,BZ/PKTGEQ)dAP,GW3S
G_)(_;9^/-9O.?V3FdE81^EM2J1OW1c-?f=2&C;Y_?Y363N1+(VWM;O>8?,+9<[[
f)R9W5dO_G]aaM)TJNPM?IaB;L(>T56I)/];_=9Hf9+.O/6MB:MT;9UC/I8_]^fa
)6R0ETXdZfG:bV._eUL@P^B)R9>4QPAG-7G6@cB=F]E/f=O8J/D_9ED&DT=.b(F+
<a,c#:7>;KHZ_S2AKI;SD.]X=gZ?W].Z1d2-:N_+^>>DAKS()9&(56Y.09_M9HGB
f:5^KIe(bac:6b^I:;\.,-AZGZDF<(Y@^4-+85/^c/><ROLK&(=G3]4-/FAAd;ca
Y)Sa:&J]+Q(2&c=.G?]fSD6)6CQ898RC_+V?U__fcTU&6WXe:<4=QVK6D]?&La8.
GHK<cAQRF4J7XIf\R<dMb?4e.f)Bd@5<DXW#7Oc<Q/-W8+KVN0SIXZA#CH^YfK->
8S22RTYBeEgRARY@]8X1<@G]]cK6B4STV3P]_B+c/U#[M6@<dfNH&C,C7_C0.])N
@7a28^-L;>aR=IM2LdW+&#La@13d^MM.])[CU?XBBbL?I6VdLX\9Qf&[78\9W1;:
4McfW)GIdCMQB(V&WPJK)6f7(PP?Xbcb-[<JSeDU,RT+.Ge_aEFX0+a0\54XZ>TE
-55+bRGTd9BU4Af4_4M<Z<0GWE]00YX#5UA<[.UNPX+.C@O&G;H^+Z^5(gg6QM0[
gb/LP-_/Y](>X6fT&ZKIWg])LUeX[<;MN9K7L_e)a<2(:2@3K:_/<B;N.df\@<LI
61&-Z3LMd:@9(6_/Be2TTT+7^?TDSRMfc8#6>B+W4K)[44>Q=YY()@^;e/QU2RCf
66Y_f2f//\7>=T77<FEGY9Z5R--2:8;@28Wc3#M9)OZ.+E&Wf&#P:</X(9K^.Xb)
cZO-f]D>S6M#K2,\]V5ATIV)b/8d7.8V;:.3fBJCeF-EP51LQM72(GM<0<7-1#NC
.=2IO7O[^#f_,1O2[VMAg1V1&X6bL5]^00=gCggX3:+-CV<9c_-W#fJH&b1_E#4Y
Gb]S9cEFOGA<<5]J4#XN):#\IAIUP&gA)Ff[Mc.JMQ&58D6eO7J6[:#:@^R7@4><
Obg:/HD(G:ODegUB7Y+KdDZJ^SB7Sa/3f2_+M?c[M)+0+.RLZN58)E4DY9P1+S,M
VY7W7^;6HP;31=YF_\>:]EQ9be]+RG;OWJ5Ic[[O/e^KW2+17K-BN6M4W2XHDD7@
gX4I+UbRS]JYRdbVEH1Ld^7SS@,@Lc)g1eVRO_WSA>&EF]Ef[51MbZW^>8/:3W<7
Z#gN:b@CN./U]EUg_JBc_1_7V]cF8VA?YH/IDP,[6PMbOFJd8]TeHGD?YXT,I#RL
dHP^MCP:aT4O9c5[0UcT^6;A4WHcX,_TA23WNO2V[aBCS;,TTb5H?dFF:bHOcKQD
C]a#131+>[V0Uc2;#L0)BIK&gZN6J-QWZPegVTDI92cS;J.]TK\=2LJ@b1=QWM]U
D&N194Z+a@0UdIKRa>bAD,97^RGd21]Vg#NC4P&BfTW#-(1C<6\;]#SUBReLD6,T
^F#GSUW_J8REeL0?HAKAaA:>?[,N2@]#1;]-&<Je,7O4,YP(DBRT[SX8QI=STB89
HCN0PgQ_a-QQ@?d2<FEN<aB:(HO_B@M_(4;c@ObZ8.>K2DR&(5f/.>_-BIE#\ZCZ
:Z<Q6EMa2&:H+1R,L0b#;[OD8BWOYKIMe,15LGOID@WX_S>:#XF1C]M7SGKB_\>I
;gIYERP=@^,UE\9SO)]fgL8IC[_,FO^=@#?-_bUBa.;;]0.]YMY+D/K(XMHX[IGF
UD5H/a:VE9_@BW46U3-&M/NHQIVN)&a)VRC/HC-FWEH,gYe;E?aa?[+;=J+05R))
GYQG^E#54C&4J]-cg6W_T/M=#KIbf_W48fM=SGES-CgD1#9g2LbX6c[QV(WB\IbB
ZO?XEXQ)Q4,0DVQbc:)O20^[]FP?\Y?Q@/]7)e3W&_VV^Q#YdRb?5:bP1U8eGQ3I
\7Y]>3QW>I86NYJ.X^eU=X@B^4ONU7LZ2Z,&P2_G>^b9OBCBLPd(D3VfM1VNI)QH
Y#f/(A)f.(X,BPP;bfMG0N[73[a7.KJ?H[<>I/?BVV:fL(Sg@#LO./>P&E41R._8
C-360B;gV,SWDaC4,/>C<6/?K-5,1J7<(B/#WK0cO;7,YF:]Xe[\-8UZfHV&d+/#
bAX2A/GG3=g]cO=W9aS9HPW4O7OIfMB;<;](KcO[H.]cZ^#&IQD6O,HQCe7+5HJN
1cc476;,Q-=7bESMWR&N-+.VBddP5dVJcgd_FY-Z.W/=f:]d?@g,S5M5UJ6P#+4_
5?B8=1a/5@^bYSg)AdO41Lga]aXV47ZJF=>gBYYXA@DA1F+AF3+D/(WXW/GORJX1
;X^b+,]_:<3N#3D_+-=H;R,ZN3c#.eaPa]TG2I<dOF8KR>-3&[D#3Yf77M21)\O@
_YJ[8FL9eI6KE;3fAV<(:&QNF4<-YG+^FPf0)V];e#,;V@<0N1eKSdQ)C:a4-JS4
9GMZ?D\b&ZZ-=D._4b0AL+O4b;06Y^;egY[0:Z4?6+H<eQX;:79]F#0bM5N.HgYB
gFN\[KMH:Yg#cY0F6[a+=?3PAJ?G:<Ia95IX4Z-WA@&-;I.1(V>V-DHa=#b:J);X
ZdgQTQ^Y>30Q3OHGQAMT4Y/:::WU)a#eR@DRP821g\VQX.PHVH1O25_9;[B_b\9Z
KKc^,3JO&&[b3eN:2bR=:XbHLZ[bMS>5YZP7U+3;QJ]fG#:FKQgQCP?FCJ\2AUA\
C8S\NeUHcG&H-ASZBHUgBQOT)-K2[e5B23OYIZ=Z[_V/CSHHP-/+,=SZ)OE08YY1
WYacDJXA@/2A5a;KT;CJYF)9&S?DFb[a5^RHQ,W>7#b/##aLYCU9RLF\#DUA-<43
[\J[SHBW7dRSZYBMU]PWT2W#,3d^,>9JM9bK+S?ONU:Qc2Cb<8C<:28Z,IH,H.@5
dIT2E(=M),OeJ(AKYNTdU;OG/eN/3-c)Jc+,VIFPID;<9;PLd4<eR34JB1P9ATTF
X+O_Z_eO[U>9ZJ<SaX;>Od=AS99b->Ra9YTY=[;b]@2YSag/R+@[@MXgQ+.>&3(I
I5f-W=,5BZ/eT;6T]J/gbC03g^33;Df-=?;N2VUX4D#CeI13Z#)=X]U\DRfc)=LX
Z[(<KfR[B39)XV&KF;6R60HH#<7O.DdTDQ+Y\c.H=-K9KCcG0DNG55;7H_QLU-TS
16EdGH^@0_M6NU3QagA_RQ56;fLQ]>CYbQC(bR]RBE;KRO4WXeWD5:O5aT0L]F3V
#AV12A(b+Jc&U?F6)E/WZOOI,.3CfJ>50D?P@aB#;HC[c@#@?/(DM?D7cC)OD.R<
]a7Z8IH2,E7&,@CC=<\][a&UX<C0J1OUW=DGJO6W8=3YXEa[RUJ.c^/3PZd&)L:0
d0M@NYc:+FcJHd-P+IJ]1/b0La0Z[8PA;U@++<^=M/+]J=525)H_^D^g+N.=EaTJ
b<>WH]Cf5e[F-K>^4W]WU(5d2ZbcUDM\<O<c^&L8,XO_XQaPVO1TS+Jg@)\IW?e>
Za.L&b:AU2BN8eOM0g^cSd,KNWLEHHd[A8&^>V@@@Ed>2A9VE0GSeI:@DT(&.DaQ
TIBQY0I>\B9ga/O>=a4;0I]K[Z;OdQJ5&9JAEXNg.SUgGa^?]TT47HY=/^I7A[_6
G]J9H>\;IW1>#LH6HYZJQ<:VIP&[8UNFI4O,[4\3+H_@>DY=6&H4@KM\/MV\C0_O
H#TQ,ZR_7?D^a?D\BFBM]^be-\_O_]ed:V/>CaV(41=0MREd[[BfKM=I=73F4_d4
#IU.I9bcdD@g,4U:e[R@dg\(\bSCA7P#76VKQ@g5,5J#_)J0<:#_9I>PM53-;#H&
8EVI8eC_=[Mc_YNRMH>^#O.O_X]FC_,e5Q,KIbBI93J;8YACKgUPTXIC3@CM]-0E
<d8MKVJ_S2MF2f/A<B8LG?.0CK?YU+3gbfI_QA)e,Y?d7fRJU>fEZ(fe^a+5g[@-
+H=PAS,JD?6E&P3GR)2fVP^6CJOS9C>6ZC&PEFgOQ(1g1W_>3_5.^AKYFXN>(dVT
4_A;2<;YdO=6Ub+K+S1ZSYH40<?G>e:^-UW0G)R&U2.L.RL7(-X,dW8d4E>K_F4_
.&b)VcK10F2A.HUDD&MgR1DOVC6Pg-f0<#0>O-c=&X[?LX+))Y8E(Q2&TG9R)7SX
RA(CBM8ZY?3339E_M]+0JY5<d0\BM@-I^&bd89YI8[BLaLSW]CZJRW0UEB3KV\@3
WA]VJe8Q/;?Z#O49P+P[,VAF)2F&[P4N.&c(c[6CgfUMO3?(@4f#Ld-K,[)3V71?
0a&dK4DJH4TQM)M5dFUT(NdD/4V=>9E,)XACb_RDU@JACO1TSZA^Y5],aJLgX]H-
DMCf,da^)0FEfW=I)CUVOFOaCaEH[@HVD0<(U[T+50We<\)EH+4JNdX/14e-O(d9
7IEKH^UO;e<F3]>(J[=Wc>Z0R-QE(U/F#D@&.85RHS)+0F/[e#EA_L\#YX.+^,)d
B(7<)&C30+O]&,aH+9[TffOR[@M=2aJF0-@cXA4I;B>>@4+UCY6081a:C(S^c2;?
@M;YD#5HgRH/V3O[[8c99CD.7W1UH[&GUd/,BUcYD4A0:88eIROV9VD4g]Y@-\M@
MCV@29DB7NfKBG,U96N8f_0YD>QD2B840GabF+3(\_3-Z\_ESfGe_e>-d?@/__a(
XZd(\NMSLCZW:9T=[SEfLTP\FK0EDN94+cM)?=cH]6G1]/;:&23LZE&gBTcU\aLP
@ULH:TRP.S=TZZ=cS(:^LD/Y&H<C]BG?L.OV7R;SJN6=gA0+:[a-Y9U)-Y2[(0NB
XK1K26^WWb#OYJUKI_X_EH3VLbSWe&^=X5-O<V@[PdCW?CIF4<X6LEM9&D7X1,1>
JB>^0<g.#HL0\W^CHXQa,H2[C>3OeKPP_fKZ]CSdVUU1?VOXD&a9),LNVaMK<3?:
^ITAJC+2b4KNLcOLIN5^fIf2443e\&Uc:Uda?<@]O3ZQ>&>I]9Ge1c63AUHgPga]
YQ9L>8TFBAYGO@e5gSc.TQRBc+XI/J9NE2c#X5Rd\6aI#,)#,Y9?Y?6+<WQ:a8LH
QM3+=DT41LAA8E/M7_7]/3EaI#1IYW_.8Tfg]1=Rbg(N55e27;XO2&-WI,PXc.R^
a^ST4Ta+cA:6g[+)PFV<4\GB6-gN\/7dAAafLb?XI308US+cFH.c:)W9WK]]>+gZ
HY9V:6d4M^SW/(<L&C?&_3af8MO0X&^H0_29V^6./2C33?#d-3]Td7WOFOW8CKN0
;32W/B2J\Tg[gW#J,Z<W96YJRL\bf/5C7;\7gP-B4#?>:GX^37T,[0g.7ed/HHTQ
9+717f-]cU[B1>PfD0<Ga9Nd^b#7V+^.1&+O(5I>GaIN_b^\61BH1:]V@)([#[;2
)c=cBUY]Q4+^5YA)4;9e+_=@W=1DUf-FP4_:=DVN-71D3_7\f.(SR.])bX7BYBG1
-2(L4<V6U,.QgHYFdC\2c?,B8+P.^_EW\cdQ8P_-55>WI9SVVPAb#J/SgPP>-59O
C;VQHaUW)&#f3FL-6_KBN/Q/aS:X;ff2#XLX2J?3;@cbP21[f;bgHS1c[S:+?2F0
N4Pd=VKNDc0ME:7aB[PG<8V@RL;9QS&EOCTeL0;@._9FHD]KS#,QCJ.WdCGa3HQW
G1IMFH_KF\BN4#8,J6J,F_>QWW.W88KU=LZ6(BfQHHQBLW)9;Kg7[;YNcB=T-PKD
ZHWJ<M=GK8fM0A@2V5]IB7QGbW&:]f/U6[bR[MJea2X+Q_,J#83S<S5H+1=Pd?5K
G=T,#[RM[]O>Cg;D5O#TG70ZR,[X4bcYJI=L5Bc-F@H]WG_]:V,\bJ&AI1N<gGU<
.-.TNBM.<\Hd^5L(R#CPSI8F\XR)Z=&-)IYM9.QaJZfG:8]ORHc<PY[CPY+F97g0
:]e8@_+)aCbL(e4+:O02)97G[L\L/+M=>ab3EJHQXGH#:138<[LOfU]c-)7TSG3L
69C^KS+[cTTSG.E;U1T:DAcH4^A>BT]DT\N>f^]R^4f&50_8,[YJ^5N3e<bb-64S
B0J4Zf,GL:9U)6@eRYK>\<DU@:NLC:33&F?4)[Q.YP>ETW+?0<=44P+NZMJ?))Vg
a@^d[T18WKWYM^P7J<@W&BYZ+:;GcVJHb(COMMTc&dO8RLXHab<K3LI?Jd85F-U;
f159VMa4H-4A,I[)HK4DKQELd[3]YcdBU=0+M;QTVN>S#RRR-bA>+R>)WQ:XZM+-
(.7L.D_WTCQ02#?DF0-I-aT[BQDQ0.<P@&R#]5XI3BBZ\([+Q#WNJ.F:-33U>+)9
0=@UV+UCK0YT,E&/G/ULC60ceZ#?dK\ebP//b65ZB/1GL^;D:61E0fPKE7V^GR_U
?-V77P+91fe\W]G^[2@4WB__0V<4Pg_.C>R5&3DR?TU:f8?G/AeA(3SZWQE[XeR)
7-/&P5_M1Y+J:@;28CVFfP2-_V?8_MeC98F^Z0<<6eQQYXE\@7=7C;+5gF[(84eJ
N+-73fQ8Y6NJ@BT+R\]]JC.KSD;N7Me1U;_,Eb]WM8E3O21F_6BTID,JV+)d5ZAN
KESC88:D:AAWM[=MB&92SDTU__#ZNb6f72@cUX[/T;.LTLK.MF8E7fBY;N#-(.02
1a0QcF:&-0SN4ff,F]I(NLYFAUU_NZ/PVX+M)@Xg6S/(\K4Ue6+g,5JeR,1,LaFJ
]_Q8C3HK/:5O:)<:2\3/)QIL]_2YVAe24OW_0)9(5C=d@-&Ye@;@\I&F-Nb@:SP+
C[K/FQFFHF&Q:a[&A=K1K=2/>D;fCP.]/Ngd,1ZFB/\f/Yg3_FTI#Uf=1[b\L;cS
fF^U/].Q4Tb/Wb.CaSRW#B[SD_LB@U5aLZP#F=g;:<MY]E?/bb-9S.=G58A+:L4G
aC<]_RM?_738:bGYP)d2#J)NO5#bHS9P8I^D4Jd]d5CG?5MLK5RcE0#G./Z<R8YN
Z1I3c<UHOL<g3-XLYQMaKTY;;7](>K_1f(1K3_RHPFVQ(-,6)9b9UA:=-EP#;V9C
FC<79#O7;T<cO_#1G=#Gba<a1(62gcQY053,O>80W;9.9YSI-.+]L12A^c@<Td,]
>Z)KXa,S4Ba.K7dU,dI9O,AAK1Pbc;cD2MKAE>8UX6N6f+0Q:5<XV^NUYELK]AFb
/06OH2B0)2dbIN&Z_;;<\>-96\FOM&6?S:Ue(0CIfHG[M^1@3QDK>@.VXcd621Ef
XTY[R=.>\f?TJD9494CM[6Cbf^?[Jbb]aO??e(OU/R5a,eNR&9;Z,5TPTI]dTTVH
[^eSe:Z1&^+&c6\QfP)2>@2dbH4f3T+CVTfB&a,NEIFZ^4,LfXZ@8^EQL=])TXWG
+PH4Ja+?).2C2JFUW+a68R5=Re(^4&MF?VP-?a_>N18C[b0:ODT9]4KdP@Z6a.^=
\._?I]+e-&W[2B/RAAOL48_]Q=RI&A)#HQ_g#@)RKfL[Ng>3D89@<C1B0.dS)3#S
EgUUBU3/(;]b3V0fcD^G<W7-[e4LU<?EI--OYX6GKPJUYdWNCMU)e+UcQ5@)/d3W
F]NPCfU<I_;d/c23/H)US)=L>McO+R-P1^_b0B]_;GV)VeJC-ZTS>EX,GgT_#]X_
@aA3aUT-6]=JI6N_eR@M,5f/:1I#IP;//ZbRf=:ASEI)D)XY(.eK902bd-3H8IR8
5?N@g03R9X7Z-KSGb1F&H0>O&dUdLM\..MCS5L8M@,KG<?W.^(>1C59(T=L\YY)F
>JR?:4]#HgDfH,.P:/[HRAA#4<(OH7[6a?>EM49ZHY-:5R:@E?B.<Z+\U8&;E1XD
SVBKJOMH[NM_A=XMLZEY5(LI&_-2\9&ZOEd4CP;dANY4YUT+DaF)&MT\#>(D2FBg
,BPX2#X@eFKXPQPQf-FBF+[1-)4&L)/P1.b#\W.+c_9PKGcH722)2.g+A]E(a)b&
=?f8VfH]\N/Cg,1(WIb6[[J1Ng+R#5Vb(a+^5+M8S\WQfI^RMA@6AQ)a?>1GR.=)
e_QfOAEP#g&.WQa7YT1>408M&EgGF+SI<7W7(BFTC8-60G?3Vd/f3P3fgZgc_EaT
.BHU&S=Q@gPM_D8D/g4aCJS[.6-WX+756?WGW58Ra6;&?.^&B=F9O7N6;3L4+1>Y
@MJIEM?/:HJ)1DbOCO;J5I<Z=@YBUGGWV>cYSUXJ<(F2d;cA++?;CgC0ZZcd:#3b
>(FF[(9^5AMQ+U)(?f8PBQ?D<5]4CU?&QO7^XHcM<A651FJ)DY7R4#NgMT7GScEM
@/bXJQSfF^0&Qb+,HeK?,?FeCIF724I=:2=>EUEc+65cJ9]6\+9b^?S(8VEJ_V>S
HM9](.#A5=cB,8_+[JQ:-8X-=;S6b(f]8Hg+_)BK8/SS5Y@O?H.2X9@&?.b]cDA1
3V7d>HWCJQ/W>28P)[Tg>3BY7eR)/09A0[JC_=[DN5+=7?:.;:SRI-PW+5\E,d0<
a1P?&gGEbbMFO-5394d:4-SgRce5(KH4bR-[-&P](_T>(POf=d]7MR6GA#0JOQ,^
D31TQ>X4F.SU,C>6cSS#T@+,L,T^T^Y9)Q+Y9;&FN-VF\8+RW(TeJ?;>>80-cS)P
#I?c\=ND_WB;.LcP2XIaQ=)&MJ,bO&2>65(FX[dL73VOXSGB-L13)O5bQTWDb^ZO
(BVP66@GCBC^HI+P]cKY80Z/TD\P-fI2=I]g9M4#P@Q=7()<f?)3[3@=S0;\Be)+
J_>1R5<O@A8e;=@(#cCOd@AW9)B3J>VDHP?&Id996,/5H/C:6+]BQCaG+R]NJTL,
D?b92X>e(Y2?_?S9SVUHScZ:)GEKI]HV1N(6Y1C42PFL9WeNNBLNR7([3O1We&X6
7DGQD=R<J<U#DV,9-1DPbD1::cLJ#XQ[WN[3\AEB,ad#cFP1]#]EfS7F\I9(+.[Z
-=e5:8D7MdYdMb)/GOcHRFUB1JD8CG_=#M.?5KI5e^RU^a3;T);I#S+[:^#cE-U2
dg,=)L1\VAI^0&U2O?AA9^@^4S2bebfH(D>QTHcJ-2#4BUba8)dBX]+)@YLN6J/T
0Ab5Y>9c\@<&.IH)a=gbP/:e_Ef#VBRO9#?B[,#E###K,<?O-QcF/geI6/Of0D(C
dU=(F_.917OATJN0DfYZ\?F03N0+LCc>QW5BEN6S69LdRJH+Da4P4;5@1R[(0dV\
19+L/?#^d;.#b7Y0VJ[L2V4(;^=JK8I\YM[_DXYKLR94G8+Oa#C\#BK1.4T;)LfB
[O7NP2SG(49U92+-N;e#LMYP-CGYLUaU+L4I?F=UXb.)Id/cE5a@C?W^GM7@DeVM
MIOJ>R^FP@e1^U&<e5Y.JU?O(b26TVdbE1W_a-GPf+M)+6BMOMX5-U]+/#M_-SR5
#Lc;bTOG0,.6J:&dW#]OaeU,;-.&^])Ub0RUVa1-B@T/A)NZCDKNeH_D@_[3[+QK
5RKJ=+KKK36(LJUL-9YQ[((,P@V@K3@-F/>.[FD8Qd\^@c?BT,aOHU8BV:WN^,Y0
CO\52,2fS179T,KF47b_HT<9G>9]7Q]F(Q<.Y(XWHZ\?)Yd,/XXg[NW><J,QZWIM
)L9a@-,2-b2O2AXLX1D_d;HSP,67<0\A.N>UQTJ.F-_WV6M(fIS3DOed88-:4S,C
4-)g=X9,VD0GF2;E6W6P>:cf[Y]H<@RE,M)>ecf&77CK[CJ(B-e0W?)B&;U.1E+e
[BX[MfeO(MIY=M24UTYd\A93Y2=3e(E?TYgI#;)GM?_(;Be(OB#X+?1Y>gA2<d8C
05EQ6,fD>N[79PH&6D\D?N8T>)1e()(U[]-?.&A.[_S15[W@X6b(9.AG/@;aH7FS
>UKaaT\6MD[)4\78cd3eRE;E5==:VQ&4DI>>]7=9^UBc(4RICH9_:JSG_?+7R@Ab
=G_&\fXfG<e79#ZVDfa)f9TY]T3@JB?e5T9ROb2[CKB\TR^W)0H^E>cGH+R993D+
=K_V);b&/-KS0.CE19:]Y,0M,V6Y3@J+KQUY_I@D7g-RDaa0U]2;XUB.312e\&H?
]DG[Zaa#IW&T[HD[DHbZ(CMf5#Ibce,c>c,71D?\@X1=+/7#TN/2\MKL_H3/X.(f
,4ZGG/e\YU#>P^I),J9HF^/@IeLfa<-A\;2=FCM9?8^O:]aNVa&);PX.64T5@.VK
38I=A<,.ZK:<\\NG)dN]_:gH(L8[aOP\E@LWN#\Q_b9B_CVd0WHUQLDfG^DG\RAJ
4eN[)8EGP9+UI@X9T]OI<?4J^(G-,5(Y.A^^9YASG<6:+6F1VF@GQGVBC<25dWC-
QSTdPI;Fgge&&M+@T82U-_+/AQMKa?.3.IdJ7E[O<9ZQBd&L>F.:N;c9MYG(/)F[
AB3Q0C<&S;O6\UH\+M4WL@6#.IXGTa/0F/]&a?KQcTSSDDTENSQKNH<XO\\^I8]Q
[[2@#QS>X&P^XOTMP&8R(4Q+/EM_\]5dd2N@JL-,KXdEM(@bIRBHT:OdaXM>#1:O
JP_3V@3)c=B:122&K@>7M]&@N4BS7RXX33&)S[H,;72@_.ddUd(NB8c(7<Q1<2Ib
FTJMTQ,Y6GUAPD2YCcRMSD8_YLg;.d.]H,^NfAJ6SDbGMRJKgeJ;L);17BB)f9MT
F@#Y64B-C^X6Z4(fK@R1DH3#NIXT)K-DQ&5-cY]>;AB6b6[df:cQV@J<@@;-dR<T
(1WSF#G=@/QKV08,\GZFd9Q\/1WZ@D.P@#1YGG:QW\4(g>^H[\?JdTAR09+LIGe>
DCF2@B_?OYH3>#@)<gXQV\A#/+(]Q<FD&K]<>c9c&Y?LV.X6X5=6P.UW1^T>R(>N
8KCUe9T]Y.M@+K>6,@ZMVXE&@.(3cg)Pf2DUdT^AHY\gJIX8F>3]-e6g:b@?3Ba6
9&:gF\dPZ)HA0Ie,L[5F/@A@Tb.(Q->&+@0_+d..VW+f0/K#bb6PPQ]b0d3SWC0^
@<CeAG[QL.YcJ>9S9MZcFYSY[)X&<EI_^/:T117NEF9,4P8gK0HOTQ.)1]_QL4FS
8G-b?>D+ITd\C<#,dNfYO)S86aRe-c^^DX_bYDb=RO<F_:QJ4Z-3L9bO0.C-0AXL
@^_Te<2@2@Y]>IFNg6G8VA>a_LN43.0SY[^N&&(A?D?4YA-^3+[)<HB[;e7VT=W7
B#2PCS/M@66Z6Fbdbe;E^fd@85HDKc.[H&AEUPMD^CD.K6=ZGH1MdP_-IHQQ^T-J
@V)IC23B&I]\,HeO9Wd2^RJN<D^K@=-1;L<d<S=HUSQW;e1bE#fA&6Z==U0c:7_2
LPa2:H4Z7P&,8GGU.feYd#O\?RId^-RZ_#<[<75_;N)M#AW04MV<0]O/2.#=IK23
CVI.b)&,2ISa4;XDZ4/<W9Y,IX)]U#V?g+VKaS@K4]D7a(\bWe10eEU]HEaV<PNZ
2I-CXGK-3TF/NTDC[3EP-)9<[#[R)4;K]P\9];?SSHcE:fH(c>0d,-;,g(G\,L]?
JQ7IC:d8eMD&GUB-;#G4EE\))b4V5UN#850TF#V=fO)UcHc4e@J1E2&=<gB@;1#Z
F3QJN;=&eF&YG4(a#7_55\U5LFdO#g561H=)1/4@[J7KLJb2ZeE_Af=T>7PRfT;&
HW=EYM__,8RS+?KRS<)[eBdCTbM_D>(X&HPgdT\]E6C8BAKV70Y2W-O.\XV9FQ+J
59L<-\N5;XRN>JYGVYg)#KD7D+XX9V[_9]BI@Y+/)S:DfO4[gS:a8#HYaX&?<PH;
-5E4G])cI2<ea-/B]8N(76R/9X,D(SD+47#^,<X-d4H)2JIR[#eF4,LUIVW(.ZDY
G8+UXW]?DU1[PU):RfO;EOC34JHG8EbTU#<<9XWTQb1W.EgYRC7=C?M[C_3M@23L
DC6P/U1@(/97-;VUB;UWI8M(A=fR>g:FD@,@;DC\ATa+]R@d\BbMILAQ841?DcM3
GN-0d]+T2OO94)B_-NO70^9[a_S]N60^f>/3BA5ZIA#;U?;L)+JAF8YFV_H::>?e
GN9:43_22M1/Tf,46)MR-&Q970XQWNQNXfCH=U]O)cB#g?42b/04M04I^-F^)_W+
gIQH5V<2]b,,3LK(VN;DEe4I3:L@&I85&3Q.?.S=:>Z-:We48b;ZUEU_fg5f=[5Y
_E000DN5f7C12U)C_5^F\@eT6A+ER?;MRZDS&VR7A_DVR6Da2bC([M-:>-(3,#>e
BEJ;;J@1b3)LR3CY90X1&RPDEI7_XXaIZ8\<QS9L\V&#b5L^#>YZ[,e7(.NY9C/S
a=53H?,0G:+0T;/b#>MNQS6A&UYYUYOAcO9&(_ADT]Lg)/K-T]XSCbWECQ?WU[&W
NCVJ3JH++-=+?L;6Q,B?)Z14S3FXG@\gT0fF0LcCNgZU(C3=F)fIER8/2>DSQbBa
5KJde5C/O:bdI;b0bB@3C\dRZC;6fTaROI9?#?Xa:eL=C5I/D(S>FGXIQO]c;NM;
d-g:NV80N[O_9EdVUT4e[Hd:0E>TE+2I7KPM1S+4UZPbDS1d^6Q8PEbK<@5b1>NK
G-(^/]9U_LD=[<N&0QR._(-df9ZMf_9@XAbTN@;5CMO#<K^O8][T9DZ>-LdKK4W^
,c[4Hc&/X;F5E?U+8HfX[,Ia=8?F\2C_L0K^OBfDeIg-Q\&R1(4B=3+9gQJL1(D^
X#_HY/G+_,>[FLeJ]d,RH\&Ef<F07<9XGUcb5=BLL-BC;.5,fJc5NGX?L2GA)Y)X
V3Ff(bUg?^H4RA=ZPdB3=D_1?9/E]N/?L1TI)0^5-&+Q7f0S,g+E@3QY<8S=;)bR
&6^;:C6\0NdU,D\.+M>@1V&?0c1QJZa8>GVBYccPOFb3G33?dd6[Q_[[=(F=P@JK
_cW8KXHCa.ABV=[03QFfJZ&)6;6WI5>K>XPO>bWRJeJL;[GOXQ2=<Id5f32O?L>T
5#bbbFGRfAKLF=AA^QR1U;]A?AS0BdIV6bKbNAW(AVMUE1]0./#^\0[TFE1PbHVD
\\;H,2B?X1^f0W9)8Scg-P4[?+CO^E4A:>8O#HH0X+6OUPX5e>,FSSH72V<C\NPc
XL7QWW<HYEE[>Z_Y8QMa8,4YO/UObXQPfU92\94=NPGT#WQV):bcT84FBCZ^OCMN
XZPZ9@,D&fW5+J<a0MQ/8TL?OVc7b]f4-FPKMX7Xa2;9VbY?D1I4AV;(22.)8@X&
@:7&][Y9_YWDfPX8beBcMbW\1?EL2\I.IVW-&5;(LXWV?4XaaBId?HZO^XNN/d?c
R#3>NI0EgCg(e-Q5T_?C/cdCD<45T-C)d/<GI-Lc0Oa\e2QB+#@VFZ_c^aEC2LGC
RcfSb.d&GFHOfC4JWA\O8PWP6bCWTSNZ@)5,bBcSb]d90(KA(IOf^4L10HAW.<..
eA8?5?0AS.2WD;@(_H1DAV3fcUbNfZO;;Y2<:E#eTDb#L+#ce\KZBX^R0_dR6T7Y
V^C96E8fAL?1QHG__#(GUYCLNJADaH=?<aE1Df?]6C+@OMF+;b1QMb6?UPe#-0;6
NY1H#8G/2\,W<H7cc^C+b4D\+>Gf2-675=.^a25>U6TB:C6ZO&/1=ZDf+aI3U-KI
ZM=BVQF8,=OZ#IL,FAdb>#A5Y9423P2g@dRGK7S0EDZ#?/XJ[g(4d4:H2.Y2J@dV
IU4+Wf?WDa/&QGLBC-QY4(OO4B(<9LTPW+JdM>6:(\NS>-D2\/&T5V[<JQ&-L0DT
0&R/RPUAA^04N&/>ZQI@)D\FD)7US:/\0T>HLeA9g[G\g4<>L_b;3E62GPd:O\b^
I/YZ+BB-Y[,AN6DC(:O,UTC?T-E)YZMFebNPEZKYC2Pd>WfJ+@2FPHe?Z0\7/,08
J0TX97YG=(fUOS:]PVWFMF.QV\;V9OU:3>LF9)F@VK&JW,+]U]B8a17N=c.)@^3B
^A,WHS85VRGU[I:\P_^fNd3=:(VK7HE,NM#)MB(6H.8_C<;4Ze<<6GO.e<fcOG_d
ZfJ]Y:KWX+W\e>/E:B6V8>Df7XJ9QD9WO5CG@(f:VAT.UfWPX/Ha1//,U7<ZE@5H
c5E=,a0>:5SJ3)ITRJ8Z/]@B;RTR;C0da;bC@3K8YTS0ff&SX(TNWE,B/NASE3Ea
U3NM=)P0c\.LTDFZfKO835KfP-Ib&W)0I9/)3KG2B#R<QUJX0>E99;NaJJGT:RL)
XT)C^E^?NK/78_[V)GdIRBC-E:_f-1>F^X#C]F_Y,L:B0(M#NaA:AgJ-L)SMGegN
1[<aT.gQ+9Z-E<Eb-9.S(-Og99]>4Zg<D15QUZUVP8&2&@5Q;EHU<(.0-A(Id33Y
E@-0+V/\=3>I/JD9bQS[3g?1NZe4[@5CV.-YG^Z>:,([S1HaK[[TLg]PJRLQ?gZ2
ae?U+f1N>AP)Ieb,EC=-Ma90Q>W@,&.PN5Uf,E:O4cF,aC<c^NXTGHP#e66KKDb:
\JC]BMN;@=VGK&#DYaGX6G2:](D;,(S+dMdbL[8+WBJC>f]\d;GYCS0P,+,A)#=R
fW[FNE?,<6Z[720,<04#?6gSG1PdeD_8_&;bSc9(F<N2cYJVM+3=&5XG7@AISA74
4H#DZME^e&QVF1FD4KD\7a>S4Nd0Z#RIaXPUF9(SNZaT&NbC>BK]aK&/C5KL3]5X
(1_2dC_KGQ/@YLKQDb)9\C)5&M),9)V/+b@B/L8)d_B)8V.KXRAa[a2\-L9WA=AQ
/C@7Z0YWa()B)EBgB[=+&K8d1]b5:R>K&Z,8YA,UfSHB8cN6K;cJgc]/]KLG(M[a
8H#,H1ONIH\dH&[\?UIW)fHb^=\VZPb@Kc;8LJ:a^8ea@KNG+L9LT@<UQ-2a&-Bf
a2Y?THe8\HPUKEY(Xce/)X8)O+<-D1a@a0,N9.--3T8Y(S);_B_64Qe5AU#X[YY[
0JJF8#T5Yf9cIR9E;G-+8FR2F.HL4KJRTU9LD&M=3ST+96LRRHCJP6&Q87.c1-Yf
d43580D9>KDeK7PSeZc9dFG0]4b=>bE\HP-g<1V)]0XLC_?6a6B2GFGB]YY]^dO&
-e#2&HO1>f<>FI^NSGeT)L]U:88eW=YMD^?YF<U5GeM4aBXP[dd>JPEIAa0H#:IU
E+[5,D2N;PAdGPOb;dP11+3RF8/\3a;;/1G1eeL2J9FS8f85KfM-(g.:BRJbTWVf
4=cK6b]VgON2)FZE?77A]/1X@f/9JB)@/OXA+2E)))/Gc_L?2_HRMF)2,0+(:IK3
)XK6@,<J.#G=22VE/^WJZ]O;BJ^ARb(.INY2TE;2b\XMfN<AV\7O3-<GUT7UXF8X
O#LBCdSeBAb;J@fSJPDNOR>\eOBUTa3eM<]b<b3:Pa?Jc\.4&<K\)Xb_/\^c+7_E
eb(0+,cXGXMQ-CfbIE/f#@>4EY<.N6O@a)<R(\/5eZ<N4,IO^=44X=J7:,;4_.JH
U2a:4.9]C7>D,LW7&-]?e;-dZUc.CSg+HVgYQ68Y5OR,,^?I])\>#W,Q97+11DSG
J+&<e/BXP)7Q1#1UcWe;R/^3&=&SRa@8=0_ICSUg67P.0LfATbTbX<Z?PCWF(_CH
)3^.26-ET4f)VR50U&)N_JLCQA=+16@-fZN>c71fNVK41[4D2(<]^.1e)X])G,,X
PV<T3OJS?>/\<WK,LXC7-gBfaWVPJ&(g3N[a=b6Z]d?OUT<E1bID92F^>e076Z6T
4[@1#_O1b_88A/&8D9Y#E[?8#1=.(K19fC<c<AF.C4&BKM:F\^L+BHN,G45[J=B#
G,[^Mg4F,a0SBeGE_b[A(.<=G:M5X41-ZFH59A7@J5e=).)D27QG1DEfc&_<#7>U
TfMg^=(a^B\MDQ=P,EgRKBK?6.Q&;(U<ORQ9@U/;Hc]]^e],9]=B50,,/C(88>JD
1B(;=IF_]:?+4QFQ(B=J>)gZL0#<J#^@S#V<&KO828U?:(f;?_95=+1B[,6R/aAg
U2(2ELgAO0bdBE@>L.IQ@Ib_#UP\W)_U(R6PLf@=)DL<A08<<.QHE\:C#RD(eI#U
&I&74_gPM#W;+c0B^7DdV[G:c(6B,F=MVg=TD?CQ+gU,&/V#S7:U=8R^8NRTGY&I
@.NU4+SI#&0a.J2eNe[KM4RCcK/]1C&:bL\Q@R]]#C]2D4B:R&/Ob15?Mb]-/:9T
1bOV7EA7\S8NV_DNHH52VDO(M0^1:0-6XZWBG2GNHYY?==J-WQ==Ma66@=EG15_;
KJB@YB6/?Ja;+17O5fV[[X._M2,e=A6f]\7K__f?[>0:^;DSMC)25#TTNF#c5ceI
g=TP)92>eX1:5DH_;Y:M_63Ue7-ZP/H#ECVfDIHF=^7Z2&?8\gfc9XY?R3V-/+d;
fQ-K\PfPeK#:7?Vf^LGJI)9OH:O1:\^?T&=g_^KdP89;J1E,S=+<]3I_BU>(LH3M
Z>Z=_#-N:bKE#X]B)HFJa>()WF#Z9_Hdc_K&fU30aEJ:L(6,>bd:SN:&Ce696FBU
[>F]7Qe4H75Y:ZAZ&SA).cSaPQW8J<@E7;W&P#g1>T:73C-<@a4^XSU#\2eK4C-9
T?TZ\3K=92\7DE@?UUMMXf5-e)YC;T;O?5A-(@JDR-_@@YTO@e8F]e,XH&F/V56=
XM6b1GHP=\g;S/e_\AW,[daCE3c>5;/[M,XR@2&GUfbP;@(V@Fa@Fa[T;2>,UL7T
W@MM^,;F^?UU?)C]XFDSNW4P)O&aH-EDFOeW/F]_/6;WWM5?MQQDfN6[FYAV-MQN
K5bA:)M<_+AW.YSg;J9A(7VVY+3+MM;.Med0.f30Ga3N?K:E+-D8=d3_H_&/6G;E
E6f]ZdEg2@:<\94=_U[C>L;ZD-?YX>-&BU_R72HgW@D16Y/\4_1bWW>XSeVa7;<7
c8?e9B?e+C,1JV+U/P&1O<E[&^NMYbY1LHA^OQ]8-3.VJW5VI-fVMOdD190-C2)2
Ca+1]0J=J+7>M30>,771;3GFPf?SKM+C2;Q8/.MZQ=K2<^fPfL-29I-HL/[DPS#b
U]41&aJ6OJOT_I?#),P;MCIXg;6.f02&--(dK\EgBX-BY6LBb-)P:;RFYB=S#Ec\
G0FIS@K>-?+Zc(ZB_RBR;JG4=OHUQD/G;G5EgSG6,XP;eZSM]6LGB.ZYVRB#G9_M
ENN=0R50;JK9L+=d?M4?FW8\6[?^eJ8=+.EOCQNcLd6QBOTGOTTg/CCfdFC<=N/3
Ed+DT3Z;a.V6bd[V1<f^_IAZQ4:L4XYTZ?JTA:4TXM\?1?TU;]@f]aH,>IGCfN&A
0K;:2-H8V&2_#ZI[WAY_6-AcXA846^9WL=)@3O:fGY]GS^B[,1GeB]EVT7UbSR<+
RTO_>5DU<_JUA]2S.TJ.,&Xd?GJe[U.S)a?E-BcFPD9&GHVK#@BWEF;aO@I90#6)
7(7U2&I&NV?&YF<=ZWV[.MEC+a-@)^e6gAf-EEXbB7gYEdYd2MUTfA;CZ@=YF3Y9
@OHF1d_^1BLONP)<[)B4+f<_BNb;[:eX)G<]&?B22?Z9[_HQ60fVV60+5(7J.MO[
(8HCJX2b\\c:>Pg(UC&:b3?a8de8+@_&Z^bWUNJ^-8:0:4L9@&8HeUaIE[KTX#:e
LCXPDN/[bTOF8W]QfTAN0fKF(;75+^bQ;_D1RUCB&[AR-DI=)?V[/+0KTWNeRWD]
6ZADAYN\H,M&.bd&S@bO>6B2#EH<5cTYAU33E[4c\KZS4\>@ee0#7<6WNKb&:?E-
^16McI&T/R6,0XXbeO46RPBbW+^ZNZS(_c5TNcf+8Y5?06.&EW-D[.(=I=Nbg^+c
M\FL)NE+gY<R)>W(C@F&>1;R)\QTU@S;U2Ygc(9T7T1K9N7(K?L)IC;ZYU@C.]H5
FbNDg^=OY2)841(]9DeQ,?E^Eb6<4L.1UO6QA??TF>\Y-cZ#8)J@V(Q^.8Z(?+W<
=3K4Y.NI>Z#6cG@OdKX#UKd8<@FMO#M=7Z885ac@CV>J(FX,JL\]a&X9dZDP[[LD
TTaTa4M?C2\--@ddW(67^Q[(+e<L)Jf[_U/XWZLQ[-0]RU\#];,IO44_RBA^e/U;
Y:\a:+MBK92LZ-7O+V<>gK7&G[)WDb8dD4U(#+c\H:#@?1d@XYI-f0a@MFI0G.E9
=_8b8>]S9N[bcQ_G\O#bC#+VKWHBbLBIN_b<4P2U2;>)-J>eIDe_?4>L#BF1bQ3Y
CZ=0-HOR2G7aDKa-S-I\4Q&>@cO4;(>0/YQPIUHR+1EECb23-4FG6\R&]RGR:;E;
bdGaK]DM9H8O44=5f]&M=[VROM9[e5F>8IUOCFB(?<UK=N]9JBA4\cbFQ5@-M_98
OBBLcJ2X;9\5;J79Y3>>Yd#3LINKeUZT7TQGG]4WPG.MIgY\Cg)[(YdTQ,=Db,cg
#6I_1<#\<L7IBS<aJg,)Sa]gL?6X;P_M+U-d+=)O>I7^E5TF49ddbIQ1:#7F8bdN
-+R\7,6N.=W9=[=R?@d>Kf.g:DTOdE4;d=]Z<MD@c;A9<_]=:(Zbf()WPb39&ITH
-K#QL4C-,8NSCg767?,P\VQ6Z8\W(PgdP3I1Fg?/e9gK42>^Ke,@=Red2=fO>F^T
O1(Q=&DOGQ4[-FXMb\aFLf#0X<+4gd7cWDB@RE]X74_7ZaPL(1G)+ZVCUKJE7FGT
:fg2[LK,g7#0SJMIed9)IBg@O[)f4^I8+W@WD5aHM>4bD-2L]Ne/0:HJ?7]VeF#a
C9Y(aVcREg5N-CQ8[\C7J[Y1?R0_I43.#\6)@IYG.XNDUH:Z>_e<XM_8DJU.T3O4
N/9<ANBCSdN@S4W[O55+UML4<f,8H2IUTL-6C=C@#4[3Q_DQgG_CL:\6/\G@^I8d
d0T(F?1]e@dP(M[N<VU0DNU;]f7b:@b/+QYXR\WI(L&aE>W5NdB\ABX=/DU74_b+
aDVM?F_VO6\==AAI<H@8#3BY?.ccFc/gReMP6gY4/8HC/36EHIRAd\>?<Y8<[P>0
bZf9=AOUVL[+&+\EM97)Q9D_39SK&^?Z<I>gL]5H/,I]S5ZA\1:6/ZD[B\I&WLW?
DAd<<;OQWC#dWT_V?T?GE]-Ye<?B(Z5)D,WG^-W/bJ4f1U2.;)FD8AL;4#D-Zd7U
U&Hd\#8R(#edfW#P36)&D(5I#7aM5M<FO(-A(\S]SfFK^V.\LVC.#g]QcXN8/L63
a\=OV0;6V=<28T.V-<;f(O3_[&aKI01(bW0gK?HXRE&^[b^_#R</2:Nd1&RF3YA/
ZVR=)?:EQ#>B@g:f9_c)-&&c/.D]],<X=WCS>P#6I>_1?E(:2=A\OQO,.-X46&)+
Y5EGTfP#6?)&\\Oc1&@KZ/e8AgKb&3YYNcMfP--KZW,:eJI5-PT+Mg0^H;?TD:)M
7)gW(HMa3LEIEDKOQfN>:1F:-dSX]bbf9/6EX2][D#UFQHTTKH=/C-gFVAfF;B]^
PF7Y+#f<Ie2]d)O]8NEIK5/JfGdd/F<I^D+M)B+<O(YT,?G#e<T5Q>S/=WM33P/R
11e6Y5JE57V8JU,IaH>@0d/\IH2fL&X(QQR=T,+HS>.]d()DDHP2ID0)-dMTC1)@
f\1E:G[L[b1>LZH8dEO_3TR4+A_5<]?)8f[>c0\?]0LRFC:O??fdFM#QFX)1,UF-
Xc9Q-5,4Kb=HbPP<0BeCM?QG4]+<34Wf+WP:c6.O>RH8YK6IM366[f]B/K19G#EZ
UF]:H&VRWQ_1@@7(N.8+PH+(S)R7.J^3?G8UV?Dg_N4f^VZRfb2bY?/1e:b8PN31
a)[D.;d)2YJVJE5SQN+S_(IVGX@LSd/J/D7)XJL94<DSg02YP3.c@:WP?#Z^>)O>
/>5.7U7\2[A[[58bL<6<HHO&_2dJ=?).,HdAFg(dP5EZa+OPTN<R_)&N-OM]5O]]
S?X8=S(+#>.V#74VX7b6(SKB\11(\P(<_]Vb(RP,-R/EZ3#AK<d,J;GYfRZ5K295
S;7d+]XagF[U1gKJS?NCUeK9&F=eg&,]&_K5WLb:WB9dKEO)<gfb<G.:bb@;765<
X2a2^G7C6OJG,X::a___EN;=4Pf+7(b+_;]7Z39/E+Lf6.&1b^O9:YQ1c==O5]W6
:=X:B7<#F[E_Ug@f\A55&N4c9]C,^fb-TUfSFP0G;EMYXX_4cLdH6-PgZ+gY5>fS
7B]SfD=.Q2VPG<Og2BO/c=I\LT9+H8Q/UaJ7b#FBL^0Yfe)?b>7+U0PHBOV_BR1C
[MQCg#A_)8668)Dc070W.Q6:N-G;H>VH>Jcdb7IeMVG;-FA)<c2JbG>Z-218R28_
49X5MFTD7QPgI;9P[Z5(Q.@0)cLR/&2JfEe4YGY&,-IBcHdVDD^)D(6IID3N:/S^
?>TcRHZUa50F]/@4D?#Ng[5>_<+UA>G4PN8,#aWb#D#WSG/B8S_J\;ZP8<\&W2#[
FLCKZ=+HgB/M,fD&^8THL0XO#H7\-P.J4;TZB5\<[TVVH4W0LK(7)0?[0Ga?([D>
ddOA\#.2Ba01Be[R_1814>,6;4,fOaQSbN-P&@CH<;Q55GTH1eI9]-HEZ]IRP].G
B9+)TY]D8.,fNGbL?]11087R:,O-_b3J/JKTZ7G@eS-b422+G3O#ZU<8?M23=SNb
H9XBR&FU9@PVG-g)Y>E[?I3SCUfBUTU<fc)QYLPW#;6:A9Sacb,FH<M:GA/^)B8Z
^PS12A3(CFf1O&C+V_C#aAgMK;5F-ER(Z_\L1+F&1;78WO:[/@]g-J^H;YUfL5^\
@cT0O/5cBSJ+-TN+g5[W#b,2M3QXKL\&cOP(g+aW3K3#^R>;Q&JA7F21=^V\N<OM
^_E_&>cg&W+F=X1HZDXH9a:;1SRUO0=DE0R6_X#UVKIQ^F9KCg796KNQI_J:0RCM
K[+HT&H7f8(A?9I7#W>d8OERfW//=?F96b8=(dL(fXDeQ=CcQI6cF^G3F8OJ=3CW
2DL_8D_a,5W8ge)E+6GKIH3>?JEZR,FgH92RTZ6ZZ1f]P7;>5Q?e26>-=3>((;?E
IaBNJdMOKE<TRgUdO&?e-X7Sc8B2&1;A#2T_+/(882FB[X86KVb-d,Z0=;MfCGO8
RX]dPWC/0f9WH+]USQg#Fa;6]IFb]O@G0+B_3/V4#\SP;ebf#2\TZ5N&(:We;_2d
f8>>;J:?\7;0gUPX1?5)9/QfW;Tcd0FIcB.Y6ZC+&g@<;.K9_IETgBK6;>E_Z_YJ
Y\f8:=\D6QL;6W#4H]Y-I[=gNJ)XgQ21T3BfD4T+,/.?22MZZ[Ye-U:^U69GL-eM
5d.?B#:9#[J,e5OT4ZbB\A@dG-L80ZD@dSMT/H9+B)\:.@-S+@X>(FG?;ED;Z#^+
.VGd^g16bH2M1Cf@J+^L</53HLBWYDd6Z>4CP]b4-Ef1\/bHc1aAJ(_]ZFQ,Pc/7
8^[=69SRNIaJQ3J]:2&@V08H0R2UZ>PAQ\.e??DI6OURgAR(/NH@+RX>2Wd,/@5&
eAd,Q4/<VPAf2b89g6JG0O_0\bVTN4\YLOIS]X4<8TLRL;C0aCgB<VME(BZ?N?)7
gV81+^TRK9_+.#a+UD]<[6R)f5=Qg6IYVS]Q7;<HRWZ1PEONTN4T<fAeL4:A=Ag#
^[3L-.[)Q&4Xc#I4e9A_c^Q,.AT6@/8;W?]];UVNVM>?dOO-4&Y<?AP6Ra;SPZ[^
^<9#+H+Ld_#f2&PD^O^AffT,AGHE6NMR5b02:Y.T-=@))d&D8KE;RJ7]]G6bdS&c
PN<g?aW&LRN6/=;)U1cU;[XRCRFU>2fPSVNQ)#a&\cTP[SgeUX^Ab9N;_#U+eR4O
\Ca\CZ_2>KC8N[-4VXd;A9d5WbADVaVQ0X+KS=54I4F?SYJBK\9L\gZQX_.?H(9g
(b9\(a8gX0C3SbDN?/10;/0822D#(<NJ@HY6]>F;E?&Va,FNfW_^a3_#51X2F[TG
]_8;R-17_V@OR/1PY3(4ga^WE#?>BICMY[^1)KL]8L(/B.7JJ;&c9NS[9,6#ZE2V
-CCdR4U=RVPB;R3^YE-17O=&DO;DefCHe0>>DK#cUO7R0;dS7]:K,R;3;@f/N/XC
Q#[g)FH#9<=R9EEV33E\VO1cZ9@(-_E_a]BcAR0dBdY3^E^Z<DJHc;c3J-9g_X5N
<)D8C&5a_UP=F74Ka/_TOQ,ZJ9H(ZJH-/K^3b,-X,bSa?1aEO4=^A3Ue;K/VA[aL
W.N-1(5f6UB]+O8/+V/BOJQBC;0_dF4I.86H>?X<+0Ad1;M7WC_BG1&R-@?3:]9I
QMTK4,66U^4/T2-F(JW?[C[JKWFe-:3OXb<f6>[3QMP7QZ:&X?\>HZ5a^&EedMCQ
ce&):a0I.5W7.L@KL44+PS>Z2U,_5WR&DJ23?@cMFK.H\2D)XC?cCf&;a?X-79ZC
@c8:=Z?E14PSYY+0Q6VXOA&XZY&(J@X4P^Tf>gTBBN:2U4Z?O73P5/W-=B\Ef9,,
f(^35LE7b:Ra[?X0ce3_/KbJ+\NCcR.#8#7LO9\PPF7c+^.)7eA=-+)a.KZC,J.+
E_S(gc?+3ZfRGJg/\BaG4-M.C@Ad\1G.323D#O-=MO6B3.N0&aX?&JbDM4J9U]2/
EU.?UaGDR+1I.P3/)3;.^g9+Y=AMFB:/9+D<;cELXC9b==Q9UVb0V1A_(V##_(RQ
3IT28QC+,<DL@WOgK>OaYE#N))WL(>3O9NB?L+bed884cNI;GY\]K5EM@YLPDU3G
cQ&DH?fUQV8IQ61e8cY_>GJ4>O>/73#3#&YZE&&N]JH5^@a@eLL/YO=HeP+d#aHD
H<e8_8_V_U]S^a.I6JL,HH[A=7JMX=0eA&:K8\:Y&V[8<_E[dWd)d&^6<@b8N3K]
O&P:P6,=RKEDU+>B&QX,:TA&?H\JGgOQ?S+5K/C3[EVc.Y:LecUC6aSeMZf;2O&/
_MOc/#Z2028>G8^SK9B@=Jd4g72LcQ_A#N<[:#_XT_#HFA&>JW,:T3+X1]fC0?AG
3Y^C,bPCSPV__Q1,P>BfA-.K@VcC?1B0#TGUV#<47EeSS^4aB?()Ia25#;-d2Q0e
d>G)W6:[M30+#^12V&@G_R-9[19M0@W]TCF@M;<#N,GIOcF(.]CbGV<V=OJ-X>/g
&STC[A-8-4>7V(CgD1HYZPY/.,&.[AUN\DF&457g6^R;X2_F9+0H3-#/+GEMf??c
HO=J42^6W,&Y=2?#+A=dOB8_/RO)+(V0+KXcgK^5BH3\JP80RS+We?&#9/<->TEP
XT<=IJ-Y<W/)<2XL?\JZ0DgTI]&[4F53JDRD,D^,=XL1L+=&^;=8eJV56C]<76?;
A3LI?S_=T76M@a(B+6a3bc8(FW9/(d[#61LX7?V\I);AT5FI\QDE<,[D\A)[P8CN
gJdP7\(LW42K/@7_L,LdJ+e0b_F_AT515,WWg1]Y=)D8_C@MS_LJ@3?FaO@TN9X^
7f(6VY)567];KeS(<94_Tb6H5B6/ZdM<,K,Yb\KPV7b;NI?E=#]V5HBJC4>5Bbe^
J+:82#bY,b@F;Hd5LdFbN8B.Z-2G)#+9PU?&#,0NGL?WfW)P+0XHY4e@4-Fd,Ya<
;5W<][X?#T9&TaB/()?0g@,dNOf,OQ7dC8Sb4)Ia-g3D4-9+)OEM9@BHC8U+.eS]
bHW,a6LUUQE;Ug\2/S,+X(W]G:&d?.5HT>)[/D5RG,R3U\0Rd-#)#NL(E_ePH[3H
db^B635^R4?<UGFdb)2Y65-H8]TH^H5KF5/-7C_HeJKM&BeNHVQ6F.5DSf<=Eed[
6R22+[Y]I)1),9FS)Gb(?.WBH3H\/3K3R?9]<SIVD1<[-A2>PRDIOX?D^Eb-a.MI
0.f:0OR7==EHT:dVMLA:-bY+dBaBE],F=0X4JC4a/+XU33)/#K)QCXWY2g7Z>KZO
Y(,Z^:PRED:8V]:4M]AS_dSMaZed;4.0C5JH2BJ5a\57.-R-AE)&B@-cN/,DQ@,&
QKFE\KCN@RQddRG4WAI>(dXSVJR7=N[^Z445b]SUd7bK,Q[H@9[/E=T7>K:YP#7O
NV8fWRd-Ec3WL<Df=<CHYAdQKWf+EfLTUNP+;JBV\=A5P8ERY_065]=8K@M6P0,K
DE;O[)eDWf_SH<S>_>4&(RJHWbU4>D/75EBY95[>7UJ53XSZQMc@D,,aAEDUF[<#
VTFDd;LUcgL-]BPGdLLd?^=;CJ>bU(H4/Q<[60^,/<(/:EQ-d69O-A=AP775f5SK
4R?6]^7(J]ED)L@VW]Y9CgFMZ8?^<R35E&(18Ne=/W2+AW4EM&Caa(<eB:VH\SQ9
W])cA[1DMH5M5^5:=bP3SaD_=d2WXJG#.#K?.R,#-#::-1,OgHc\aRKdI)^O7<=[
5ca[ASVY4+\A>a)3BP@)QRg0W-J#Q)dU)-T^IE)D8](]APX5F+OW0#7MAF\&E4-;
6CGBaJ7F.GIR;&E/X0/JGeUP,-,];):6.W6HaUO9O(AB?4fQ8#cU2(,^1a0W=([A
9YfP6MPUc+]a3EJd7&P5GJ)(+dHF,YW&gJB/6RACd?ID6d/S>C3eX53-8.<ScZKR
^ER_?YMc:+&.0;#GW1(=:U2c6-E?MN<M;;5:RK^7.J@+/KS[>8DDT.)>=,(2^e=2
5PD.Z]gF./)Z?14A].QNH>I/E.:<d/UM\5&62>DY^F&W6Z3RbACP6V97K2FKZ0<]
&X=gJ&SagR9e1S5K(E+L?D>7Y)M,4/TDB16VMV]2J,C3Q).L/@]@/>=80L<H^09C
CRT6>adQ/DFgOd7[?E^;,4@Q4^L@:@KQA0TT_K[7TVA0X:JG-RYE[Y8JW#3c&B&H
30E+()9O&H\WR2<fF,e5)BW>^^(U\@(CN6J.c+f,SLU=Z[2MO9,H.&NcT3gR]+)&
gPef^FEHLMEN2\cSJ6Ca=\9K\e&LUHY->MA4WSQbJ\@4<33.60_C#5+D;Uf?<-^c
.#@,Y]7I?I6WRPM,>>6Y>_Z:e;c0S1c<D822_.If+570-)UOf/HfW;ZO.I&SFGDK
fTSfB/aB\@2A6;9P4cN^4S+H/\\P:K)M.e^.MW(bK1dN,R:7Qe@KM2JH(.LU-.]-
PI_C6D9QO/1fG=<47;+[Sf3Z=eFL>E+:[+A?8](H@,8.5A8GIDc5V8fDfY6d;Z-I
KAPH/b];-73X^eS4=JdWWTd2WX[1R&VfLH<#44L1H/K/Gd<EWed44/SfLZ<KCD[+
/TPe?<9MPC#A5B5T_^2.+_3IXBafY)FK94Y7DA#W?+g.a5A0=(9B4E\R4e(gK_4<
64?Q7BJ>KPN=/2J3JL^;8#;P6P,#>SdFGXA6(H,1V\Pb)Rc[3@X0<,NVf@NI_g+1
Y[AAS\?D?/fd)Mb\1gJ8bA(RQa/U&;XR+\-.?aWRMfQGNC\.>G:40?RF<6-cMP)e
U);UT,YR^>?WTKcB/&\^5G)9_e0459=bf[fE\JG]@2Q+WTT=T?7dPXIN,5U9A2YG
&,PP_Rbg,E_^fBQ5OcO)9C[;.SI<ZRbF>=S\#8KcAgMI1\)?J;H[S2e<C\5PA-3\
6f//6O0)3TTPdNFBX)/7WOCH,dBH#c_J?1J=B5;@SBdG\FCae@Q-IY=e2&RXdBdS
>M3HfD8ROfOd<H#;UV+>2d=Q()BeQB&UMRBY^9QJ;FZJ6.S:9gKK1YD7XN23&&<>
6G],A_KAQ5[;.1.6>VD@#N@507GYc4IeU;d7\T&Pfcd8T\.DW_<(--TU6MB^\KXP
1d4IHHWR+4EW0T-=O5SQNV9/616\/)03\;E.,H+B7R.dD97HP-cEUHX:)Z3ff0G+
L(.XHWI,+2?0KgO_HAc6g>\eSW6C#;HZ0)[QgIO[T?IF7PLEUVHB)6_,7^(V^;#,
-=0<1^Wb1Y(8V89G35\\#,5LYRU3&(HN9eeP4R#^7EED8Mgf6#O;95WJGc+8)^Y+
(P8BFX=R\0Q<2b.OO-gWT6CFWLY]A2OP/eT/PHERIDWHD,a>(+GT?c2/5GIS5?LW
07AE:]Q.IF5d,Dda/+fQ>D<6<HNa1:We9X3+<f[D_f+E#68_\0dCK[<]RH7_#6B(
2BV1]&U+7:\S_J,b)f#=6,7<SW(\)3=DB3f6+07I,dN0]=DT;_NNT3<aRXJ=@R/;
c9CGgSc[O9G1KN)/<(-.V;1C_eZ-P@IPQ1>FH>,6EOZ/S&M4@\F&@1@<FT(=b<C;
1BN2\JAR\-U\#@==c1-O:4RN=MA/>=E,@4B@[D\I1R1g?dB;d0BbR6L,e:T9#Z\3
YJESDPe(QGDd8YD9#Qg9S<ACMKQXgUD6#Rd.gID;9L;A3,-G,XRgIF_2.?#H+(-_
/7PY)>>4J/?QRY].[,V?&Ma&f89Z95dg.2dQ<6/^e:C,-9OCe-:P_@UK_KQIXa;L
;:b@,H:dGA&@ccf,?.^+^=U3]J(eaX@^-.d4ZNJ_B-VU5VQI_5[/VP0J[GNNQAVH
W=<7gFb?[/T+&M,Y\/E/9F)gNL8):0L:6P8FCbbLB/RXEQ?.U6,daE2?&[[ELTQ=
dR65_Z3T3-af(Oc<<OM=@_fKdWe04N:IfOc_NZ6B>f<6e7NP#-YO3P[DD2c4;:-c
5_NQBUM]H\gE7H,:g)(ISIZE4@8DMF>HZZYK8V^9D^#5BM2,?e4?FVc9I-37Ee]g
+=G2VC#_GSVGF9\PEdN46V#??=L?)fH82<W.K):XWVSJK>;f<UK6Q??U05O/JQMY
]^N6aXW0..P<PF)O=B3=L5JCc[^FBPSVZ57a#?Q73/L6&IH_\@BK_Wf[g=\DCUUJ
[QSK3P6#a\#XHf37gZ,[2H+MQ_+--JY^E4<#_Qf?HO6b/)5-L<Z.QDAQg[dgO=T7
;F;=K3)RD2+fJS?(;@(&2cR0E+O\J@/0PG9R.<;eR7SEHb/?>H9ag3-:e1bW>L^[
;M4aI1DT,<QZGPR@-8O[/9+K-)bO/?.0NA8&XJK,:,]cI-Z(6A5cD+>[X/.&RWTP
@K)L7Q.Td]Oa>XO:0+D(BLGe:cX=[++6#>N\F=D.JX4><B]R/>KYZ(fW.c&6+)ag
5QYf+Z<Sd>MVdgLZ02[@<Z)S3<17#5Uf<Y@CT,XgV<0<PfNTR;+QR59026.;7VC<
+3Q3MK-eRMC[>]cO1U4e&G<IENWf3/A^,M0ZAD/Hd8d(MHT_PEJ#&N#gM50GIEf5
+;?d.c;LA,R0_N4bD),40)1Rd\>CV8^TG[BbQIKHC&4>HHX.HdMSH;@\27[,fV9_
#a9N(Dc6E_Tf_KR:-5&[-)XZ4EAJT7>^WL_SaW9W98]0.RD+<R9SZa+Z:YbSeS2)
S=_2\XVH.c_[@/W_S:FfPG\MaWbI.OH2TCAcQ=;;aT_Gfa2O11cS&&N5HCJK;W6@
4^LW.QeE@PB/.YA4a,R@JW)X]ba45VCfE13^,2<ZK:gLfIb4MO1I0VA3HAA3N[-V
Je9a8)W9efAEXJYO:VDb^DE(R+c/)KfZ);g<WTNcK,KEI4[ZK<&XM&EQDMN;[c+0
-1d]4SPKOOL46W@X<65MLJ]LMFD\bTL=LY14E>>.14K(eU,(IN::-(1DHAI+.C6A
bdU)/9WTJa?DAVM3GBQ]AQ)N.#Qg[]GOc-I#:</[PN)Y48#@\FM63bb9N;IHVY\-
./\_1ID=gANN_FWW<SKe8<R9aCd.Lde:=fIU.3FE^2SCa-X)^(G0[T;S9Y+O:CSD
UGK_#eSHKT;XAga0@P8,@Wdg<.2)C?V7LB&Xf4SGI?5T692DS#QN3aIXNLIOD&\;
D1/134B?+W_cWbV83M3^eTSCV49H1CPD,gbceBJ1:<9>L8,HSV4H@b3@H?GC>HG(
SVfYFY/,=Sb\FUFb?KB.fOO@2PD_12>:Wa]e<ZZ,,T:&97-16)_IFA(+23DTAaJJ
.2_O9:bCf<Eb2SS@)P8[590R(]\cLGMV=gS)[EM_<d)-2X_eg,\W_=NKC^WB^LT>
d(:;D.c?^\]8/E3&GH_V4gHbV/6+;-SW9U5=OMVU0&U/<SNALMIDJAJ&:Q#.@3a>
_9AbE<a7(:6&,8HAGUF=7.cDXP>T2]][Bb]a^9<\Z@?\7=W(YgOd0JO-gQ68/BHW
^(QE=2@\<e:U+@&0d9;8F<<XQ7(dU,[AA127>7:<M]Y_;(:a&-[fTA.CJKQaLdVH
7T=^JO2e<QPGg@)DWL2RCUf3&XdCda5LTN<JHLUJ\#]g51@BeX(BB/07P><5?GC/
X1LI\2-XO.K1H_VDYPT)NFT@7>GF)5L2-L04#IVc6ZP-.O30Ya>SZ;S_K(#,OWfH
\9YLR@1-_KNMT3Te&aHFHb[(N@?KF3V[dSK_TPI1RK8T/(&/HF]12&:_)2gOE.5,
;QWH.c+PE@N\J[L9BK87ee&UVL-9e11V4f(>D^MH:O;O:geb)S+<;c?86/DbW+ce
#a4ffLTZZ8BK3L;5BOTS,&e:A0bGM3Y[^Y>)6b)JG\PJfJCfVU,COeg5Pa9;:GVF
&afH=#INK^]4#gZQ2#:4Y534),F.c2\7_/CMT(5-S/Z9bD&DXfT0L#O+W-3gbdLF
[Q6_KT?3IQ@G)4W#K4X92\e\ZTYd7;.0]bT-ESLC[KOY27&B.O/b1RE8&VNY+(Jg
_f97H2b.[I=^b)SV5aW66D#T^E\2)CXM)4Hc_dLAfabdE#(:,;Q-JP>/PQf.DG,L
LQV8>_GOV8]2Oa/T8PTBMbYC<.Pd+TaQQdYGUe<8OFCD<g[_#(PH5B\CHf64b3S<
eOEWOGBC50/->JA[T1T;WM6]72DTT>@K2F]d&_6Z1RM#S<28H9[@>FXbK8cf)OMU
N:B)N,?VNY,H4+#.VN^;K(DO>HG#3<FWLH&1]]DASC4.1P;PU@0;).?_9LGD9eeU
.YAPSZb@YUC\Z\LP5U6\OJY3B\QEB;1XY-^dC9D\MK:F4DPTD+AWQ]MF>4?G?/KW
AaA5K(N#2G=VG_.LMB+4UOGT1UaY#U5,UfXUZMg5.1Y+f.Cd5WRFbOFY?_0aGdIY
fN&SC=V28LB456\L#T6[Z:e@c?CBHJZ^IL_;R:)IYCU7@7#g<F<M_R?X.WC-5V,;
9<FeH:@1KeG-6Vc)_X,WQB[YDJ[6^I^fG@=E<fTWNAHF(7@)M7[PEHe19YQEC.4)
VH3U.d,e)H25@8g>S>:gL;WccVSI8eXQ^Tc3IMP6W:J#?(5E8c:+,N]K,J.)[a[[
^cAI^f3aLTIJ^E).&M]I/&[?/8a.@UFOO-JSJ>C(GW=A8[@-cb-S4B\TVfRcD,<N
7MggSR:^?acA+_2cI+K_3E84J@7T830I9=1A2,_S0X04N@:)QJN.c/C2:LW>/@eM
L>;QGba<6SXTN@9<[D<Y,(69-@>,NP7.QdHT::f7?@g>46bdGS^J<Z)Z7=1Q[&>8
@67Vf^#Y#0Ybb2/GQUWNMHQf@\W9U]G;f,8d)#Ye5dSQ8K208P<U0(aV?,K0d7IN
+D#&c.R(d\#+R<T;7:IfBH]6>UWLSf::OT<9Q@e\-?V/I&(B/[=&684Y?;9d+8]S
B3T+C;^&a1TA>T_0?6O:>DZO0RB<]IA@7HA+Z&a,J7OabC(4P-&OK=UNe[_,B16c
-IO],cNC9JY)6HI#>DVD][X\0Ha#/5W/#5(XgWbFU3:Y&E+_H^^TIBOU/fTETD^e
Y)(TAS]3(0>:LACNXA[Z[#e?GRN\+DH95-9B_O&+L^c?7Q?.HA3+J3N=L.=471?R
^PO>G#AP\S(Yc:d?3SF66NMM^>Ug9FZK]I9:>X#A]TZ@D(RMWd1LUFA0UG()I;P0
1e62>4@3<&H&W5(UdY/#A_H[C]^WL=1=B)[O)\DB:XIg.ACB]..?<+#[20B]K3;S
7B##L)T,8Z&_B_GB&@gR::]5N,AGXFT@gR,]4HJ&X/.D202MD#(:&T)e8OPYg;=L
\B?KG+-JB<6@5?,[9[;a=.L7KJHG[I7Ag0&S1P#;F@47AO:=6Ied-d8]GIQcO;-K
b=Y;c;CWU/AU@LS1Y&[N8dW#C7=VcLR?F.@MOUU_g(DJ^JS;9@^G?7F0#d,PJM^G
:@AI9(4ECH.B#f.=5]Rc1MP>g--&/HI8FO-2HZGO?aPRFbcb^DO]b9?4(a]EL8Ca
^MEFTdT-W#SU1^Y?HQ4OG>K3?^]QQfHaa,Q6^)G7d\VggdT^::R^0X9498/RcN=T
=8;^<-)g+WJfLRS]@Kc#TfIG5\_JQI=?-YJT1E8_gL:9a_Cf;RB;D\fcR)M7aAB?
;N+3=ARXSU0Sa5e9&54fLDfH4Wb17E^5M/NU^IK++>7D1P3?]RQg;5),F&WJKPaW
NA^PHJ]c4Q^6<48,>FKPDGc<8/_gO#a=MD_18631#+C72^6:^;1UY8DFWIgG6<FK
g&.eXOILE]GQLS;+bX_?0_\586dUT7&ZR29S0D?L(fE/XXGPC86D;KAMe_PO9IC6
690d7(]M_^AF(0P3P(WIfF@^=.0;C=LH]&65/B\J86QI7d(eCSCUD./IBU24EBRH
O0UN_L7,AX&?0(N\6AFOKW.EL1]]0I0(H(#RbO&UOFOW/:KJB0ScE;_9IIeD^B:B
e9BQ_MBSCP30+U>FgOB4=H_PAM^[\d^IO-D]3YLe19&Q2ZB,K_9P2d#<OA7DZQ3+
/_>O(TE.LHcQ,b)V(0g5M&]<::6S&B7F]8&Z\6Y<-]^U8bHAX;<M]g#=5OH>Ld=4
Y[HK.3&1g6BcZE>ZHebHZb#[I3>[@UA\FVcd;MI_+b-^)44QD(^=cFT6#L63Z^S1
CUD&Y2W9a?AT9_fX#(e(KEU[WWedGUK#EgaSUL/(L;CX_6bE,:P.Z(-(gUK>]M)B
E:0]SDM.IZF:cQ-6DP,1S6R:A;eXDY3;TE7QedJcd.A@G#I:30b.ccUZ,VDD#UVC
AggF4XD&:B.LeEZE^48HL/\^JQ]ZY\N<-#G-HS?>K.Ig:B6)JL<aZdJ:;KW8g=Ue
OT1HPQ[#3TC8aU,_I/KK=(d<;A,ZHNfPN0_fIIFAO2-DbL<O0Q4fY5DBI#7M#&DZ
/HLSXa(_<?6Q8D6)5(#PR9g4:b^W7(/[gM4YB4@1/Dg,8F:,;0KC>?dTCQc_+R?L
B0b7]4OR>L.0K#W&cD+;B>\XLeVS?\/DQZ2aD6PU5>V_8GNE)VdC4J)0#G1_+03I
:0(,+8Iad#c_\YDBS3R_AF>7HcL7Y>;,CXEJP]a1Y)QH<S8RaS7aK/2\;Pf?+Y1T
aB^IJMOHd(CG;,T(2]-+\AfKYdeR[S==c=_3C;/XE2_F]\/b&e\>[ME:MA08EBUG
Qb6/Zdag4R<W-YLI5=TJOD3+<75=fK@G2Z,BYGHga>>?;:#WKYV<QGMWXKgaJK,R
;(#;c;^I6\La#M4Q[[X5D(<E<>B\T7:OC7YI8-9>N8dcGFQCK\YJ&KG,PS[3Xdg#
L6:XTO&A/)+TO]-I?_c4N6g2&g[NE)_:015LePBb,L3;O=8#+8#89W;V#I9T._ZJ
Z7@^F+35-G0@=&PX.<cC#0C@S=N5)RO1d66\CWWfg]UE=2U]A,&DE:HaYc;RDRg;
-(PA]KA91<B8Ba2:gcdL6V=1\H0+C?S>a^(E;GOY/3BB@EADEJZ5L:V2T,V=_e_M
9-SZVX=,eYIC;I2/69(fD:Y#C>27BKUGT^beUf>(/EWWG=[,9>4cV6UgCa+&[:3,
a3.Mf1QYGa9L;TEa[C-7)B3^1D_L+B86e_BcceEHUCG3;C^eQ;R5C\YZ:.Zea(4:
BUX+KXLa@^K^&CTMU#RKURWLHUbIZbd(^8[MRQN3O;G=GUEUM_a)dC/5@W(TLI+8
GUJ7f)K0)>R3C,=),Vb^>Z#e7@Qg1BfGI[HSM27@@H[G__1[739Y#gb3.3S4,1a8
_LBC>Q,9MeG<:c.W5LPL1(OA2#B(R1PY8ICc7[ATXKVT,F\CP.(]-.O]dcRTB6)1
NQ1&XJ):?e[2=3&)K[I^FZ1&51^0-JDJ=TA)HX5MO6Y3c&6N@-B.^1+-7[5JL/3f
McE->]O<8e:V@2MbI(;L)F5eLeM3OZR<L_&V=\[DT0Qb75f25NQSF08[PVac.0EK
PW;G3:X:HI=CcXK[>9bbZ.,g5BJYWILc=SJ[</TcUAe1b,d,C0Q>PZ+JDP6aa;GY
DB)aE?Be-\5M,A.0C/S0K-)d\ZR^SbI+.Y]6CZIGaI-><65S+RNY8V&9#)YY>MeO
2[;7OS:]FWC05a0Gc22SX\EOaO=<2:+BeB.b6e&7PO45:9Cda7\4KQd3ADH;/[C6
[:W4NS?[O4X4Q1gOC(\W+NA<K<\1IC#7D:_QbeJG03d;0M#EU/N;\-Q,L71L;BFI
DEUXa&d+H1H4PC4caG3U(=e_]YL1T9IcB58698e5/Z2ecMT,IZL//(1/=TTf9e9)
)WUG5P<-cU.FF=\R466S-aAC81CFa;O1YO#HVFXK?1;E.(#f).@5)SWVa0)bK&5F
bHDL4U@ac_][4@JHN8,K:+?+G@,09J0[4NL0]/^X4R;MZL,(a@bcg>\@]ARBA<PU
9&=g3RV?E[1MT?c.^a[c<@WRJ2].JfH3dB/aO@1OE8JJR&;IO^FO67,X59V^X:O7
K@6FaR\G-+)5L;;L;2W@MGQ==_/JOLg5BV>^Q2MZ.a6-H/?Z&V^[9D?Q.7CQ<:7(
Q1A2d1AE-Q2WQH^5TcVE:-U_&]VPbQV,&9=<b,X#M5KB#9[,f\47SL;PD@(50G53
cN=8\&cI3O4VMd?UZK@a?.8#&4eBf[6C_N2:.DYYc2[fQC33TRKQS#QG55c16.2:
9:gTaFS?dKH)W5K.WPCWd?b#FU;d;M,d84\L<04)9OB[DJ.dEPXHVM0g1=Tc,#M2
d[(E,=HK\U[&@cE-JD=Y.Y5O2CB=dU:I_9]YLg;56VGaZG_O#D]G^C\0,#7AJgJH
1@,]1EKGRH6IAZ<N.J=Nc7#bMP](fBS7O#Lg_5FA3:QcQ3)#\KLc,cH5d7JG+>#S
[3JA_6XMPB+AGb)L4/+Ke#cJ0-HKJ0ge4=;b8LSEdK5>O79^4WU:Q95#MXPUIH#K
bIA/4=Q8K/e]MHTcRQ]Q&N#S=)8-V.#eHa]bJC@@:&L5E[T;CE<]Q[dfVIR:&(>Y
1UYEBOaFG\)49T(OX]5d6+41#Y69O=aUV<SPRdNU<&5LKC_301#;24C..RfPPcPe
5(Y;>Qf\Y743/FIWH8,2dgYRGC5@&#C6IS<,H:.;L(FMV?:#?\#?9,B7.YVJc[Q-
62RJ-FPY1@f2#1NbX0&bIMeC+_X5+(C-LADXg]7?U,TB-83F=LV@7R<YRIV:T<^3
ZCNE(GHXI1H@>:GX5/NL@d7g:P\:UO+:ee-&XF9Rb,2T[VBSa>HKcBZWH#=W/)aY
cF15W2642[I_YOb-B+0T^E<Z)O2WCBP7]<ABWIV[AeAg3T1V=]081S@\fT9(<S^N
1#WeGEVb8AIPe=)S\Q7.#5N3LKBJ?d-YDFPJOR)7Be]7M,g@\<ATR@Y2;9.R-P=&
EaU9I-d/b;60X5T.RN7GL).GV]F:GAPA<T+A/GTL^9&=cD4^&cNdR16Y7.C)eT;G
3KD1COU[R#MM1:-GI3e63I=3c/MUT+MDecU(YI?UP=JX>?H8<fB1TN^Bf8T1&/:D
FgZBdeg(14GPc7-@@>I?N^#B=340.C>>ZPAgJ(/@]a?Ef2URTJ.2)(B>HQBB=&U<
2Z@AV9^2Q?K#_H_NH4Z(&U1eb5RU4HVSC&EZCNJ4IMY&gQQ4D6H<3f(Wb^_NP#YY
44KeMI<4IC0I2X#=Tc2Q)>TQ-+_,LdAQV4NW>6J^YgI7MKAgg;QMD2)@:Y,P3a6E
T#IC+00_G?X8DKS)\-c?aDAReOK8RG/?61_Vf4F2)^93/SVf1MgGQ&XH^L\;WK7,
][T\SdOBfbfA]M^a(IZG45=>?.VE0d_VbAD1BOe9D-EKa@&S-<UH@6GY=.NSDR&N
W]O8c)+:KcV^=aJO?#V=N#<[SG6,gRfBPW&U;DT2)CFZ/SOTPL#[a/QU+14L5c._
DE5E>Z&-cUKDc[fGbPG]6,S)Q?WTLf,/</9(R@cT03(6L<D1HcbK)XT5e4KBeG4+
>?7+B83HAcS=\B<TEB[1JNE5>4Y4V.a2\:LacF+XdE)1_E=K8\[f+\:7@W+CJP:O
/26BH/Z@_57)LSQW502DVC=:cN=-#)#c+X&AT@\+Xd/9G;\1Q6P.ba6bJgDB<-)f
Z5PXX\&c^B/&&@3L<AR@BgZ[GFOeKf\A@J.^G#4Jb0)OG/F8+0V7<\F?BQ=U:F-S
EONL4K6fFLB.VRBFKWL/8XCXD/c7BEL-CR)GeM[P,d>RX6&K0.XbcYVV61YDbO^(
WNDgI)IgOLS&DANT,a.J2b^3QCQ5A_<HDO-/6^K=J.(U8K<2I;aWeZL6e+>YVR:_
\UN?H1@I/9BCMWe-7dKD/&CF4L:-CW2>N.Fd[bP9UH>NE\Q2];faBJX+QNGWOcVZ
a[\dd2:S:C)T70]&MS[Q0]JX:]GVAg,):b2)OK1E(67([@K.1U34[43GgS0Z7EUH
UNNDYO&8Db1E)LSYSF5WKG0cM)f?\5TPJTH^S&ZWZ23SKZB?I&S0g6eg?<fH6TG=
RSNL/L_;7f3eZM&0,NK#3e46NGAO[JfA,SQF7U&CHUG/]cCF0T^B1J@U_,93-+3?
cB0^?eJ>ZU<SWK[C2VJ/93O@M89\WVaP;Q1-cE(K+d5&+C6f_)8([<0?<RdIQ+J(
XQ9QGaGZPVZOB)CYU_8I?(&R27-Qb+I\Z?3RTL/)6P#OMB>\/2_1>R>[LDQ\C-aB
b04/H9cD1->-N_.T3;<\Y:]ST8\UJY<42@DJLY#Uc<3.+/IY1Rc&W,VYC@dT8LUC
L,-XTP70OJa934K=T:#G4K>I]gF_N+[XL@EM8+5(BP#9+G<C.P,@))>8VfQe:HaI
8CL9,U]VGISS:A[.M4?1dJD5=N&+;5WW10gT,^1d]<_5+4-MDH6]AASD[e[=.fbU
2XGQ/a(Vf#-UUKR;e]RU8TS(-SU1Pb+If9g&.&a?2b9N&@4]O>&H=4F(/04cCXA\
W8RTdZMQ2OfB&SEf8V?(DA^+^F3#Bb[7,Rc8SR&f/:Tb/#[DOBHb]ce--CA#g=(I
CHVG-CHGg@5e+g&1e<XNQ@.f>8SX(;SN;06e@_agJ)^(cM\bV,1<8(1D>19RF[G2
[fVX;&-W:J#f;RP0NAb1S70NW6;&)_@BB/Ug&++9b_&@W(-C:6_]YDM/)(=Y<S&N
X05d7;SX5ECb\VI_O2]CH4/AKTHYROeVT&+J8.)+?)59<VXJeV35X(_&4ARHY\<I
=];F(N->5#XX.RE?OIXA#4d5<:/;]_)@POQ01O&eO#I(/f=d.#B-eFT^]W:e=7?g
B.V=POUF-W9TgA95FM(SaLR0J)->79aHdeJc\=WJdVQ[1cY]b\K4EGVC)-42R?0<
R##,].ZQFdB4FL\1+Xg?XS:QL6dPL@G7=;bg7+Y_-I+0/[AKRIN/AML\)]ZSTBV7
/Ud^C\V6&TN>=)cPXT:FMeIDB6\e>7#?2e33ccD9>KFLITSJXa6[2\=-^D#[_.cN
#&LUQV<V:Qge3fF^YA(IJA2I@bYD8UCDU]G\,[5@Db6dMBS#A5C.Y/5D14fI,R[;
,/defRR#\?\f1b_EP4_FC+\c34?Va3H,]3:9IQdAP]+JO]\OGfP[GQNC&CJ^X9b\
^[.A9gS_4:VWDe?>:GTJS?IQ4_fWfR(H2Q7>?]VQN4)@f>(>dVB&g:()QO&-B5EB
Jf:@7<]D+)I-?2Y1IRU7@9/<@4\ID,M/2DB)<TK4Ag5+PP>b^3=GE:UcIXJ-a6#T
Sf3K&YSH1ADSbRJ+4D1JQ<@_,YI^6XPC/,de,F1-40I(^K>S7[K;acb-,/KYcbG1
LKa/]8MW#Sab(D2e.>_b_.g#&B&LR9WY,UdIX+>_d12.gD9LJ=7=_)fMA/NE..Td
DLYX3&P+MN=1K/_CK;dRL&)gMMS#RDZA@1=]b4YL^LD4^+7&V2&c8Z8C>?aVFXO<
?#f_CY-S\&<F71J=8F\Nc+H\bR8;Qad#KM;L+PCSAOOfN#S\-\cM,_G8PaWL+7Mg
>=e\).;:GFdaTMBO?1@E_d=IWWa/D5b?C&S(=:=H<1_N9YB@ZU=6X(_5N.<S\_LM
dU]690#5DeaPgL27Rg0g5Y\KPJ8JX#eC]X,JJTN#FeBT57THff8N1()FBg]G)LQ)
FZ9T1YEWFfHWD_(fS70(ZdNf[@?8+cfE1S3]<;DVf](E@[M<C+VTYF@6BPN^IX-W
&9144L87[I]NB9<b,cJ>;BTBd)(^E0F=DE;PBI;GcQYQ#KJO2<9R1+-N\\):^&,H
U+@6RaIS;[R^-d@6F0OO]N78DYQPd,0^IIX(7Q;CgfGH?3Bb-)7e_&:^d@I[<;^b
:0OMe6]c:CSCTJ56)A(]JE1+C_NJ4R-1a6)DY]+-L0:A1N5DeJTPe)]-<&0P^^Cc
^^dR6ga;8\g&IV5M;G/TJS=)(Mf+Jc#I;ZPU1dgGN&CgeRHH42(<C^gRgNM#.2U=
A+\\e&P(L?D_X-d^2:<N5(J58;]6O?CF5K8Q1aL1>E>\;)Ld/]#UF=>:7=2Sad-E
;&#5B\9/1c+XXJ_QNHW-A<W^7:Fg:+V8]eR&O@Y0?TW:.Bb54&=,9JQO<<Y:3e6e
U^[0:#[RL6N5@_eK2XO,H^[W/^>YWYa1=ON_:gZTI@G7f_2fWBeI&-Oa@bd.NKFe
QdW[CWK[FfKX_P.JR(RQ,T-2OP#d<RDJ1:>Q6_#W7O?9e-PEeC5e<4M]).d;;B]U
16SV8aPc<f&,N7TEgYX2_G0CA<ETgUB05^+\_>;;1^8@<-QZL.?4WF2fZ^&C6VEZ
=De_XU]NW)O>1-RH4I/gV\#O^.:Y3:NcE.[._TXS;cL3)+Ua;U]X(/1WSE;4NI+f
&LfN[;U+Eb3+a46]85Y15UJ17MBSZ@M4SbX.IbQa1aRZ<TbSVb\;2P[9L94?F1Fb
3:78B0eQBG7ZFN/f78gY]S-g)>0&I9>=A#=O)EU5W:/Nc?GMKH=X1JfSLHEP@.HH
_Q(E.F6;D^e2fQUZ5c8&]5,SC.^dCQ8dSaF:W8e=_<Y,M3&T&BI;QbfUa6K/OF)c
NN-/MNZ=7gKUXY6Zd(I0&dRIZ3ORM-I[5QMB)XUQDXUZRKD\fF0f6O1\-L]69=3R
0[P6J8ZIf7.6Y[Z28)3MH_A[\bgLA6QN538e;f-R\5(C_4<e.f6FdCg?\?EE@68O
4V-;=1E3a<ZM,J=<G^4\@</FQe0)E[@P4Meb1C;f85KGXceYbY_24MB_bQYf=1@G
-BRM:;VbbJ.H]N3a<GKLYE#abLDg=9V+]/GUa?3-b,WY/I+H?M_^=a^c8F5cB^U-
2C<@_LDT0,JcB8QW,]9A/0f@[^GdbUaAgVTfCc,VXMeYGUS5_&A5H.V[O\H-:JD2
C.A^gK8-B,Ze:FFc5#RO4\Pa]d7](09P9X-H7)U0cCIcZ8;WU9^Ag,&<PJeT)4>B
X?Yg0C;]S]?FRe4)=C4,5F:N?C<f4/0T6HG_gZ@FUf8\YNeY_eBbI_.SLT;?/MZ\
9g\089+L:e(KIYG0+))+NP,c]JFY#,Z(d,PI.b;QdCQGF.FT#3.NMa5TK;JT7<fA
0@4QM;.8Z^;,V0KXV]O2^d759+c90L#Lg0>Je9c,3,#Y,7XEV/+;.J<<:L[V54W/
^4gJaB>5XL&R_1f_4L[X4cGFOe?.TFe;e=33-,;W(R,/Be^W>c(ca3LeNeQ&a7<Z
@BXXS)_J=aZME(4J\?>4KH?PdVg9J&IbWg@=S_U2eNV#d]7)//.O/38gWfVR&?9E
SPP8H#^##EPD-[-=g/a=Y0AJ(7Hc@Y-DIQ^7Y64Z)LN7JaG/)e&Q_/FA],7,ROJ0
,U[:/)8VEWIK>3@9E-8[@X@(f\d]\MJIN3)<agE4SB95,e15O.I-dE8RG<3G-U3S
VOE:G,8>G,F>>f2[SWNR:KKWAK&Y3RD,6BV>b)KM>4-K+f+C\VU@TL@<ZH<MaEWd
VQ_3DC)<8[Wa,GV)EKBT/Ca\_ge)7\I-]>ITXP#K-9#P6F^[L.,Y?O4F/N+025g+
e?BZSaX7L^:SD3A9:4.KYN9@V&@7FaO\#5WEFe-VRLe(M,GXe)+\\AX4gJT-,Yee
BA.3DPd-#9F4:=R\XZ8QdQ=^ATdfdZ<97G/TIWHe3QbIX\_\-)JX2/.&53;\e]K5
)?S8R=Dd9?/g<8/T7I##]Y\T4b6A^<cgYW6YC#70VK(^4P:)PJ^B.I[^()gPBL@1
([PCETVOeH9006_:WdRN/BL4L^UY(0<EFS:gbZ89YJ-V;<.0SXJRG][,DUZ5D3fa
8/.CAS3(?SR2^/>NcUY\>MZ./:JZY:&aIFY5_]8-H:.86fV&9cV&+:0^KE>>&>W/
=_^;S(L[2PK<4=XA4+UK3()9Kc,dM@#T7ZIW\g[,Ke44F=@PY&Zf^R)bPL?TOLON
?50C@.Jed3EUHI.UaE(E<0K2J8[g(A+6_)V>=4OI]La<Kc7;7R=71L>a+63M_dLR
#d:L6S<2Q<,F71:^b/@FbC-[NP9-Y>BX)2BUTG7_TMWe;f@],3,U\>[&YW2)CT\^
.)?^+N=0.5<&_)D/O>&bP@)Kdf@?/LOBHBRTC<@6g-_@f&;.)A4U26D=_g,f30.:
J3S7aAAUBM[TN3^EQIOW0#)>_CPg6&-BeUPPDa06XWM;9Pb\T(V->Ba2GBbB+&Ca
fYJ5Z^YS0.&g6;AA^fQLC=3/XW#OC&4aX(3dL1I#7^B<PCSKA->)Pf,4Q13,@#0M
OC=+G4ag2CP#\X4LH>[@1>8JaC^7CTTE1F3@_ORKUJK?_IVG^6?E(35-PX]SBDKH
B_gcY?7W6KGHd@))\J+;HWR,d^;aU6#,Aa_g^2YL3caSR;fbfX,P#64,S];HBeV5
W,,bZ@LfM#8Y3cX>,bA=fI?fP[(ZKe;[O,8ESA8?9>O^Mf7BQT.ROUb>_5FRZ/I[
:<cG.\Dc<]^)TV7#]HMdZ/M_,UD<WFY?IJ3a_dZ1#;WD#V]A8;c]+LRg(b[1]5S.
C58Z(aBM8e>3XFYN#/BF;eIg<0;/KI^G>SDg&SCE>+O0C5BgK27I(5e:BX#f\U;O
fIUF)U3N^>C0F6b-WY_>C@.PJ6^FH.[/4XL)9H:+>(WB,+Q]]CPK+aU\OaE),,O0
;9dH85YOdOB2;[\cBUQ0U(5Hbb8.72;ALQYG?cgbH,cJ24/R2bWIO#Ae?FE58CZ4
R-\(D6VcEcQ):SXKP:4/,T&S@W8d\\6-\[#TW@Pb:=D=abA7@>^?C@db(1)>6@CE
AOO37A&A=UG_W=VFWIV]:\/\aSSQQ,4B60[7T9J/Jb\0K?F;2C2XeGB_<+Y.UHaQ
\K:H[\QQ>X2HT;JY;X_L6f>9?CeHC6@#J=BUcG;\&df(K6PE)PG0\GcF=HeLR2f)
CE9GRX^S&JS,GLW\Cc(_]CM:NP[ZZM6GL<=+\I+E4be\F<B@bC,8;eA?H_Cb3:.U
PT+Q,7#QT:bD(M414^TYaU_&ff/17a?UV[,]]+_aHg8FABZ>Qg7aOd]bQ5Y:A[c_
>eH2ZRY-CYJTKY>Z24+54G[P7/1CUg;_BQ-4JNO&1L-(/Y8G<MV#/K93.P,ZMdOT
@/8\Ea(>_RcfTe[.D4OXLNCG]H?FLA[<9-&SdcIX>=BT^a[PYAU=(;476EMc2ZL#
1ZW?C1Fd;2Ya6BdF:e-DF:22:Z^#2NfPV1S+Y@R)<Ga)O,AS#FCg/5+Wa(T9;#-W
^STKd.Q>#&?UXR6>Q/MN@&,e^Gg,<)A&db5L:)^d\E9M#3PE3[>b.Q.H)TT:f;#&
N8c_IHGO@)J#Yc\4V.1VN@_GI.MH(.<+\dZXZ+QMFOZ,-a&&9Z7;,V&4YI+_gcgR
GNd31]=H9VHaHeH#9[9)8EI]_T\;^1c,9LZ)JSGaB_EWG<)f:D0DJDRP-]Vb)8bO
M?(_S_?AUd5SA:DS.X+[_8>F+C(_C<:ZIZ=/GA&b&d[<V&P:V3I+UOT#69BKZNG3
M@dRZ03RI1&IA9TJc\Na#L(bB:[6<?D4a1#RZ82fYXHGC;/[UbdMU0@:0S;_:S=5
dVWH.aWf:9B:Ib&a^?M9:Pge.=<)WLfWTV[Y6MD;KcAV5-8IBR87?g]>@Pb]E.bQ
TSMeHG,=4,SZAPMN3[6A1=?FaEXL^\QXA#aP/O)_RWBUTZ5<R-,#1O\6WYW5#NJ6
J-a,O@MAObG6<T;faY+/C<?S)K=F=MSIX9:O8B6WeXJ_P3:)ZZ[R3[a6PD=VgPfK
:2@#[=A-CO\:5<<?gGgIIRYJ+QB4YGf#&-YgeXg=5U6NE]cO/D55&5Z6VXX_^BW7
HfE0[&X_C(2af/BO>1?(6:gaTU3aYO-=?[BMP5T_1f9PX&bZ)_2:OT8eTd:@Nf2-
LTHfNY(0OKR]?MCD:7FG6DK(Z2SJZ]YXZ&_P:98W/e_]8KTAEFb:GAW>(Y8Y>+1+
dU2WQ\-fF@+W6X.]C<)aOf22+1WIQ__LaZE)=?>O_;6T0e=RcND:WG7R@H=C;@4Z
R-W8:?EBZYQ\XXO)4=2#+D2?,3D>aae><D[g.BSad6&.QDKKD:&\R@eK0BVW]OVN
-4[[bG[>>(J[VPRZ/V984?1eCV>1HbHeMOD<3<>_Q^gDA#ege@^LG1S.(IG-6J93
=T/+[\-JK](3YUA7J@^@Y_f+#NV]Wd?H3SL?VfJIF>)#.I5_B5?D?J4]#)C@_+PE
C6/,c=#3b,#EcX]Q9d=d:RY(_1,U:QJ9RHF.1,A9EfRDgaBGPK;F?N/S30#(5LZ.
a6Q3\aA(TTNMR:L+(gM1@JcH5#2C.,[1JXE15&YRU6U/0-T#d=5/QgEW2a#&W7AV
H-HOVYO9&8PE9a1gR1RFOGc/&E:6E(87?P(.:INIJdL+NN:c1J/C<J>)2fKUaB-F
4a#;^A&CKH(@:AS7@:@Ba?18QJ+N7X.J)8b6X(\AMHV/+EQ@V8KfaMC>?-&;Ng>S
#9=E=CCKVB>a]gH^Ce;9@UKQ0XV#7\eWAJNU7EdW\4URaC)]AA^g-P;?R;9CGDN8
L<fW<e_N\SbGL+:WR4,^R+M9a:@DF6<ZSDY&0@bcBb(JG#/QU12d^NQV4@)F7+Nc
1]2.#DJ:OXE^YN[eBZ^,g;I[IP8@acE(D_W<4dOX1#4P8_;O1=OTd,J)16YSEQ8T
84Z73LKD>EB(6-b(WfFO@VeQ=LeM2]U.9]9)[C>:\Tc7+bWQ7>[50T#B>VJ.eJX[
2eJ9D?@GYfGZ?0gZ[dH^@A=@M45U/_H\+23>\PO6DXLY9dPE4VYC;#2(92BUMa&M
5F[A^.b96XPbE944bfd)3J)1Gce?dQN5C9>X6W:D(>7^d\:@)5@452D@;;84GS47
,;8O-F-^BEeXUaT&23#a_(M.e/S8;bCXYPQUHT2fIIA/_:UNZgO3V&(G:27D[V:]
[2f/H;U[7E<H:O&YVTO+K?V_OF_ePJMZdf>,,\VfDS:YNBM1eNW&O/WJXP]G;[E:
?VX==-IQ3Ka\LVE@[_FO(64cAUM;SUR<XfJbGDZR>e>PPb]PL;<^ZPR,D0C;@2S.
/2^+KD:FH782RU+=JKaIR7WQd&Z])I_:5U=9GU+48?[(<(#^:V3Z\UYFAdTMBPI1
G(5]=D8VH&fGE;D#ee,C):PP.5R^E=3V-U/7V6VBdDOD.-@ILWSMZVQdL1)J.=MC
RY(YC]Y+2CV^Z<;_O1b,CdZZXCc8[PX3P9Nc96I/>XV3Q(PA0Hc.\gI#cOQITVeU
-_1d15Y,d,-LgOHL]/;fgS/e\J^K8[>cD&6U3,^@^KU5&2.?2ZeU?3B7OaDCBLc3
^QN.QEgQ#R2KeJ@[&d]Y[GN=.TMaGKCX5P1FfX4IMVZ=3&]:S^=-B2,9KFML,ffV
0H<+_F;a[@-IO(;)0#QP@Z/^-(YS&C-]VL86?X8&5#F=.FZ7++a7/5.JU78RN-PF
00PMe?U3CT9VAZTbe+&,R)H-/SH_L=C34(?]Af[d@gHVRTac;<=J4X@@H+V>,/\2
deTN)S]332XdB:SPDT\ZKF@ZEZ.^X5^\bR4<0N24)c8\/9YXCCHH,@:(S][39A^?
)V98(7c1A)J_U#:LVaW>OO<Ag66a8J3X_=7MXUM6P/QGC</3>NSF3>eQ#<4H/-I+
U+U0\bg-]JPJbg@eG[JaOF[gPe_LT.NcL3D,PdTeF];55f5ONUHQadI#Y;6H]^RE
.;GH@K7IcX/BYAaK40@&BKSX]5^N]AUAVTISgT4e1N7d[9AdTB1LC\TNS<]Z.d@A
^_-_&b]3M=,=e>/M\UE8TR=+(4,=RTe#a(WW0UD@C(,T-OM(M1LCX/NKR]PNX6Xa
KT>F;\49fL@H#GffTgcg1BK#9U@)0)M7SYg8]bKSXEHK1X3:2=bV@:\1,Y7KM5Ob
INS8L[+B9^8DV(2(I/eJI0NT3,IB+T8YM?_&CTT2(LN1_Vc.ONb81>dI?M<YRB2;
,a2@B_eT<a=E7?:_Z^2UJ(:H.F))=VA]OW),,1N14d9._#5LM^d^O>G;7N>Q][Zb
+-R3g-IANO6,1C8HeANVB^ZceO2d03aIf#BA1cY2=UBOA[#ZIN-06eN\UeK#PT<S
MCDOYW;[DNcFX)MC2F_1+F#(K7]5]M7Haff<KUD_f7WG/2gSe_B53d2,dbT3c=7>
g2&O3(XUSD1(W#LA2KYE04H>Q/1H@0X)aP_.0bDJRJ6a@P4FE-gWAcDgfP1+WRC:
W0_D(R_>T?Y?7G\SR+2N,0E3cW8RJZ91=1\;TP-_HUeb,Xd>=E5PN&fDQB>F1e>3
+[b[^fG[>.:d2>1LT.5aHC.GEeggYP6<JJ5gO@;KDJ&7)^\I4LYFF4:_3NF7V]Oa
I=0DVTHCV[&fND^?3[E3f3\X(4gHL_gPN/25?TAU7SO?O9[C(>WYdV4ZDUS2;Ka#
5>D3@#]W^Z<T1=U3T>FL(6c4QQ=(f2V2OK=+&(3X?#69V.?#5bRLF.RA++OcLgK(
[:=NQ2ED<SY=TML3@:59(??aNS8QcIX8_XLYI7D7N<1Scd#UT0NPN2O+,821)Y2I
6[#e73,]F0&Q\7(M,B,b)d;[X_.5MX<NW<AB6f&6dJ;(NDM5=E.:V=e.,)<;0c#V
G)O(]GJ5#&_-I((&C6cf:W?R-b.<:PDBC:0CaAe)_DbVND=BGb^d#G(G5;^N;X2U
ZN3d1)-YN2,WCSIYAg]V2[0R_4[a#?&[LUK:WI_Mde<ZCDP@#2dME54Pea1;;&9_
K>QR54-V(UT8B../TF8Ga-T)16gfF<^7+3>YCaBPD_/H:5)4:@QTDe-c6CcPW5U0
e021S(24e8aZ0IF93O@O[>\-(HBE,;D1e8M)XR@;,f.Ib\G)(L_.QWS#@)FZYK_2
:B/9ZcF:P>L-@3SD8OagM^A(A[7\EAE52cN\VI_5I#d#[gU:PAcSfKF.JJ<.N?XZ
K?,S+W7RQ__]7=K+];=ME<RBJ+J>adTd\8OMa86Se<Hb6[T=a.HYV6a=..6/(RIE
JOKJM\=<V(^?C0X^:EU1(ADBQ-B6@4YeHgaX58GJ(MDKO;Cg#3eRWJ<U^3C2WN]4
M@;@L#&0-=a?ab/Y_Z2c/F)gZO6]B>CF7B:\_S\,@2aB^]LO>]LKC</S(P1aNF\M
^/fB4eJSX&8F_#1?].YcgL-WCfTPdQdb^Q:gd#^3S1a.cZ)f[cP.IR?T1]a+VKT#
<NAM_._2fY2g(Zb5EE524fN1J[S>DASBc/R9/Xf=T?Lb/7[::[FS>e?aPL(38F&J
BcZNKQ39IWM&E-&E\9c7[Qg-f9b0G^.IQ3-66aAIZ5O]_:>Mf;MHOB>6EV(75G,X
VXF7;9.?[P2--J0HMS_.;#HVGEV2<I+&EAa-2LIK,Mb;6-O]BIBS\:E:W,\SJHIR
gJ-.)N+,g_>RBDH.^SR>=..:?7DX,EUa=V>:T,F03FOXg7BBCg6K).D)>Tg\W6c2
L,WT16=fMUZ7.ARMH8UKRV<?Wc:^[-X>]>eY)/19aI&O1bIY8d]MJd_/f_>;b79>
.N@]TA4TOLFXQPb\\^eV-b]?L==)fba[8^6<D8J([L:==-567)deC[1BTgW-/-FT
^80a95Z_C/(6)9&Y<\P#OC2ef,C70UdO:A8aP.=QfA(^d]S+0>(U6Z8QcN95B&d&
gL2AdPZOa5KBV)6JGN]H^G1GMf=f^^;>_0XD49SN4PP2+Y[&B+A0MSWc?gDXZ)CI
[e&dT2ZQUAeBD2A_;:URSPZ,C^Y=Q>dZ]2d1TPcO+)8Ua3)bE99SWX6QE\G(P3S\
H=CJ;@gZX#YQf6gH:T@g>K]Cg>&eLG9EL\3-PDS&+1<\)9#LAacbK><>S15KUeFQ
NWJJK=@49;A-GE6M;SO/CC?e<G3O]AR^8@5JB,3G.E;VJ]CQ/#]7QFK:-N1+dNM7
PY+bNM-U@H;3\VHSO,e8IE>dQZ0d2KB7U54.[T.,YMC[<#g&NF_V\@I]A-c3P&c?
I7b>c&V>4EM&:0]GRG4I0G.D8G37a5[,H2?B7&?,S+&?0g]EY@UEWWQ40F]8/-R<
8CH#FK]cBC+S,A<)2BSN02=T13/dP/fM&eX0WF8)DHU?KD[#^Q-:(0)]PbBg@U)O
REI-=EH#UaFXH?T1NM&A?6T5:\XD2d>1GJWC+^d.XZ2OIH,@D1cMa6=<H&_.ITG8
g25RF&8Wf([.15bgWd77SYXFYQZH9_:#=TPO7<HS&TH@ec7&DTIPV==:SPO)A?TJ
V+<g([YW3YS4-D@.-=-])9KHADI+CQ_^<]L&8f0^NN.a5_U3.X)]8;-W^1bSK8_O
;C5()5^SQ+2c,BeR1E5\(@Y(N;cC1HK:U5UG=>T9@R2GAT/]&PNG,WRZ.F4\5<RS
c,JY@WG]ga(B?Z7NQGM3Hf51CN)/^=?Ib&XDT]6W#+MQaf_LA/;4>TZ7RLYR8a7-
M):bR,@7:,W\F,O-@K100a6Hc95MSZQg>bQ[]7M=&VMYM(..2+UQPCA)C8V4&,4a
?DK?ZV>_[HLOGU<#F(\?V1d;eb]ILRfMc&A4MY=AdVG1=f#\E>>+,,^RY3;<]9E:
OI2_TOXG/O_R0:O5()b>ZG>R#N[RF:WA,=7.=,Kd<JSgD0:EeZ\A:425ZCX@@2<L
:0CRI/3Ze:25US06H&.0aL=dbN8<D\bbH>N(HQ+L.KI3OdRJY7bOOL(-=MMJLcaK
[-4[SD4Eb._5GY^-8QOS.b6-d43XTXZAM>FB4H:PLL1@3bT.-Hf(+:7<P/?](XJ?
eSg#8TL6^:89[N\,J9OHQH(7cJ?O7QbX&CZ\f,_Q-EQ7S1-?V(b/LOb(=>T7HT_5
Nd1CA]L.PB_0TC>dbWg_e\cBCb/L]Q7>DDH2B\&^FMe,;YF)FKOW87B7fK[]7J=^
N@V-].DE(_X/+(bEcgSJ8/&K/<]NV79-[(2_6[EcWC3IUZLNF=L>I)W^72UD<>-B
BRNC17VL@PRe>/KaB)@f?HO#=Ya<R@WY3Q\\W^WK1G+F/N&bCOM2NXPe\O)bdCGc
1&P@JK@0([;KG?1>/:\VXZ)Q?d+J>5e0U@7&7F?e3]/[IR:AFP&Lb2(P-\eJ]b:/
SUC^8.HZPP]WKdOabN/OM<eZX0Q+\(]S6g>S]OA^HDMHg-]-3W_Z<NX/0aM6.E98
<9HVVS36-?-X-YV=]1Nf^R8\+>Mbe::OJ.f4_bWc3NZXZKb/L#R_^,P^PbfdKR]e
KT;9.SB)M..V]]@TMS06;,TSL.D0beDM+IAK4L7#6,Tb\Z7?I78Z8X529F_B9;_d
54,6T&K?<;3,[ETN72ZKUU^0da4F;H(\X[K]J2[UY2S5?6KI_)CcE#c=dZ/9H0;/
+,7[E7/+@^DfA1c/@<+2^,(514RO\XHWI\AU/[@PR/aSX?:)STb0DWHXC5+O5@5_
)VQ<=1FGY:D(RAW,-SOd]VCRY^BSS)@NHZ]?<VHeQHT3LW9c4(L[WKV90NOVI+9d
aVS8DT]./&AWCL^I6A5U#Z&e7eCQX(X599T:VOZPPWfefN9VP^e)40XI?gcaK^gc
&700+PV0:_QX_6/I#P32B?8D=Z#Lf+MNS#I]XS^^5TLY,.6PP/++b5fZ0&?C<[<.
D\8c9a\03@;9G15ggPJ&]E95\W0?df:A(CNWUO;^=fADEgBQ\gg6DIYYIdI>SNd5
@&BPaM^035[X?<<::O>g)QG]QPRV>22=a:).WX_VB0KM?4f:Ff?a_Z#ON:3M/F.,
g2ab0.04DYN<_Y.7=ZR[&2]D0=<BO3e93e/JS.:S7,;NV(N+7:&JSOZGe)&LFF42
=8dL-1+Me.KWYV(F]D<4<P1RHgK3LRJ,8fJgeK)Sca.a[3b4OUX]\a19VBY,/SEG
W);^EgHC^RDUKTeF^e6d[F7HD8B]BK7#c52,a(YeQT04+XXbcgL=/.CHF.ZC2</F
@.c\eD8bRPR,IIH1G3-/V@D23)R:VF1Ob61B;/9ad;<(5@FK=,+G<R)AUCV>AC?8
[BV2X7_g^E>5Ge,W#E2_&fe:K5Fd)[b:1I<?:/A8(.@Ub]1&M5c/e?ND@1Z#]HZ]
52O)A_VGa4D(&A(MRTb]&YG/4\(0S^gN\/L\gIaD]0ecUUBGcAdO@?J,U##O0&^N
T43Y[@4#(eSKJW<Z36;Nb8ef+aXIUJeZ7\f?C61\f[Fc@bId,L)R4Z]OOAIC-,_X
2NMdS&N3(ZJOdGF8;-SLL,<W@:D5._e4H-/VAP0^gBb8(aO10=,=/0DZaOM1dCCM
4cUPT-DK>5g944EfV^R<Z4#U9&C92+#[1J1b^0#GP0OaM#9M0g]<B7F-:ceO9?=;
F6&<g^M5HQ4gcc:Q^g^Q^_a,YV+/RF0+]XEg3JW6[J-NAR]TG/Ld4g^X<;3O]9]F
f(\M\-g@:ED=,RdbZ#C_M0W0f=9ODG=)I0G;:XVU4.@H+G?5bWBE_aIOPDeI1&@3
@F5W9&R@4YH4RgVGZPZ#2:gFdV\=[&PSO07:dQ6]FYbQXM?)R,JaD-IZ.VR)/0,G
(C&<V0_,(SS61PUT#^fH^4_BL1UQg))LCbO?cCCI_7c_,1:6H.UdI.g;W[g7SP/a
&CRIVN^(^LcGTT;O#V[060g3ee6MIg_g4P2>J;<9CgTg2-APTDQQH]\EAD2[<PgG
I#)c54#5730(FB2(H7;E)g@@LOE&-3O3N)J5ROeYVBJ?[KCaNb\&U/8-7^<6&fU:
-9>-K;XX3WVF<>[(@MOR2[V+G+1<:?#^8Q_YaZgQKZ/4#@L?3(J?RND+/cMG)GGJ
S(0\1eEOU,JdQ)1c(2bTbD_P80QB]@-[3M)82O8WLCJbJf33f?;/)C=5</=Y9:O9
<W\>H0Y94(^4\L3:H()?G</OgCB#)=.-L,4W_RT7AQ_K[PT>ROR5;B()??.LU(]1
PdBc_c,a@YDZ&RgE&aY^eVLLDOP:M-d\J@.T[9,#S).)c-3)S()O9&B41Z]K;IC0
,(5IX+5N<abVbR\?^0Xd2M5[:R2)1K<0L0+b:UfC[LdH8f3[PNPd@bg3T??0ZdDK
N1-=^BPa3(GR9:.YOWFP[N>I5SfR_6W7Y@dL@\e>^0^@MD@?L)G0H;f_D;d#T+,1
/ZNA_3NY?LI2d=CNE7,42.56-#W_5_(D)1TUb5_Q<.R#<H&^JK3QcDPE.Lf_,ECS
7M/M(\(&Ua(E0OWB#D,U1(UQKadGOUZe314&_5XQ3@d@L0S/)f)UZ4I3P+[JbS+W
]Y=3Dc:+&fCTTc^38_LCSa)I6WFPTa,^.(bF=bIcUL-Y4H)XEEFc:BRUBc3TV.(1
H0GQ_.&L1^0AC?W9H,I,_O;+\&?(;S:81bA+Oc8@A(ZRM/H-Q]IX.5g3@TcJ<PK6
:TMbYFO4O,1]2E^MMd])5G&Z9SO,0dPb>V0@1[aZWOF(HMJDAQ6,\>EA[E[-M470
gHYZL;XeRCHb:NVBWY30GW>dTXQ_JFVIW9eNO-ZEGD@I#c_7)+=-O_)/_0TCbcE>
DOAAbd2_5;D8F[^PS@3gGL(KEG[S^&PG;9<OS^EFO9D5J6K-4&ZQA=e2>J>)]5U+
N?OGHgELHg^cW@5LF0cV&7>B)Q^?REgfL+PCS+Ac@T&4#&VF;7X8YQ#<7OZG[YP;
>gbJ;1B2J#Y&9SF<S^?4PY7O&;_K0K\gT2>,2QbXN<HL;/.1LaF>SV??d?;Y6TRd
6E;,B27Z,V?E9A(<?6(G[M/:O?+QSc;@dWU_d71[HAbf_G#H-T+19^_9aDY-JWL4
318#gT,;12&G/^@bEJPSPZSSH@]Z.W0W]^HGfEOM_:5<6J:=YGU29&&9PH_>Md0(
aD&.&[UKGaITb/:=?Qg@GWES@BdXE?WOPcX8_(+0<?\eQT#09cc@:5AC&E](RQ[c
g:SY&-+,fcL]9>e?H,--5BA)@I&<-[GS:cM@0B\eM2S/A-S,C_e7cNd.,>.=]^\]
=U&LNMZZ3A(A<JNKD?CaRHY,XKT70[O(F)cWGD@b4KHbH@>/IfHcUJ&.==#d--V,
Y9(9;?1fU\gCMB)V=-BZ4;1M(DBaFSe?7>K_..],1QX]GGG:AXV=FNOa7O5Uf7TH
09&fW\_d>e1QL+UW;a#XZKUSB@@Rc()/XVWK-K25KOMbOd\Q#83F5D^8OCa6ZF;8
@48:E?OMNF0P^2Ka3M?Zf8KGaXNA8fFLSZ7E1#0MF&J1AT:\c,AW;dB>gA:F)0QL
C91A-)S+Ye[c2OV11-</NA/Yg;Y,Ka+cP0T>;-&cO+ZYWWW4R72IR2&V@BX33DE]
aCcIC@8cN9/^16Sf:Z.HD^>bO=\XBPg2c_WEdce&04V53DDHFM;-2c1-<UMZ/aAZ
<L34<F<+f24ST\:;U7W06L+1.eG,+@;Q6HA2LV(QgaF@AX[H^=(W7L72-Y<bTU(7
IXP.(F6Z\KX[V5^WYe.P&b^H0FC&_F@)#;>GF(OFeb,Wa<8La56K4@EZW7^e>01Y
OY?N5?aSdX&;cg1/DL.gF,Xb;(7T[]5L][VLOP/]><C9M+7^g65;g^/H1OUPUbJ2
M^T7Kd[6JFT\WdF>PH2O6ZfL0&F/R^ZKT&fb@PY;-QV9CUa@&a\7B@-+/f(D9W8L
&9_SA4Hb:_?+#Bc5\TgZ#9>0?>2NM?cP.3^K]9VC<J:Sd>M1OF-a=@-Z2&&fOc3f
g\4E&KS-,B#X(U#-620(+g;Y;;7OQ15fM^TAZ1N/Y\D;aRF-=0@5B(PcYG8N3R&c
8,F9&Fe_Pf<\,,;83d4W3Y81D_:A)>2TJ9R7RMgG@FGW2bYP<7cgXW[EN9&7KM6S
&P7>^STcG,)1/T3<d.RF(J(bGa23L6LGSM_^?fU5]N>Q^&<VWg8L8:@G\B/THTCL
/AXG>L26.d.+ZJKd6cJ@R3[]d;N4)QCSSQ)=:]6P/YPS)a<X=NQ_Y-B+=UL?2\F1
^JWC\T2d?9J?Y/.<IJf4Z8,EB@56@8^AbO8cXJ\c-=Xa5+--8C.G#@WE4X)Z>_GG
E.YP+^6]J3_S>>868<(;UNZO>VS#I@IA0;=N4NcS(7\N4GJ/E2^bX\)R]^6R_&==
0eHee2]?Mg#a/fI&&N:>+&]MEN1B^gAGAbO>//0VB6T\HEIaJHT=.STcg54K;MT&
1;0FZ=?E9bNM98F]<G9_-&#5J:=dK3L^A7S,5P?PYf>HP::_]8ZZ-TY#1:2.G1aB
7P^N1Pdg[>NebOTM<g>W5QI=-f]O3Sa\.;AYJXgeAaCBQdS8IeI#0Q<+4PZ5,2H^
7IO(#=]TW.LK2J8)+82b@P>YFA0.ed=,Rd:4PI2B/:#);Bf]-dW4^/bggUJa5D?.
2Xb<1#7b>MXZ^-@]LC+[_=Oc-B0Y(9&511IRBSY[OIf6;FM<2O6[M>YCCN3eAOg&
WcTUK<B9Qa7[N3S;4IE^\GQHA<_:S_(TW0D1&97>GIE(UT<B#BcE;9IS[4ffETX<
RMLYOZBGaYO(_a^0NRW1b)R73&:0_:TC0Q\WI6?fZ8PI\cE+9N>V\=?La7,4aRX2
5NL/C&X)54af7<1NaBJX2(KHA<07S+Q9-5&>UT,<IV^E.\9X[I^D:G\dI+#a;#BG
]C^/;UI:QWL-M,+LY.XPBN=/).#g=:C^6X4G[^?Zb+]@aXE/I+5)7E)EBK]a<VLC
67M\[U_5W3G(3UeF=B456V+Vc)--BaH<F7C[TRceGNH6f\M9_FMB<5O/TRYYX7aG
-1/,1O,/?+N9PC&Y:YTNG-&ID12S^?Z:TTZSX25QYO/<Ra8-9HXU]\0OZGP3ST1-
Za?<P:\SL0RQ]4aG8L\ES5E+,2KGL5;:9D[;Ke.c984+YYUQ]A_&],dc=P4FXMUV
&O\4^MT#9ZBI7:AE(]^Y/c4ZG___2,K#Sa8;eBHJ;>>X+I>e-3I^MRJML86@O[fP
DY[S8aSA5//55+^110bTX/4fg>e@ZY@^YL9/]Y?8&,bgW0)1A6@9PGF:[=3I4/&@
MAa(6I]U_O+4<VHNP\#9(]=GEH5.AaD?QWC/<A+Dg82=d?;PW(+2W0(f/O]OG:TK
[_ISAa9D.-Ea=E?bU-7&/C]FG6f<;eZEV/0UD7;MEZ#MSRJ5>(_Y1<7cE2VW2V=J
MPJ>e,59IX,;DOPLYBX9S#OQT+.^I7XK2F652M&BWA3FA@ANS)B+5NT0fZO/d?eU
;=^gTa=;_A9SD@E:5X.B3OZ9f4A,1?g)/0>OD8cHDCW]NZ/gFeIe[#b0L98MOegP
LO]]4e7()ba6ZbO_<(Q/^Zd/.+]1[_@A>)JT8OO,N,#CL<9@_S8#=>1bEdJMNAe>
8.2V#D&3GbU@gT5?c+4MS#1.)BNY&/-eKFG,SW<UG_DODA1E4SSEGO0URa^N]VU&
L4J_D.PP#GN7@)DA/,(\8:d+c8OMdF&eOgba.<Y.7K8VYIYFK(P_PMA:ADUdRGF0
[O&/5O.Z+\N+9@?.RVM&9SfM#5R8-W&@,cDC=)b\27^A27OFB>\3(dgGA25=Q9SE
3YIW#6>(8e]\;/IU=]MT#)N?),)H9E/BLf5>a(PHcI.+K85^5T7g8H05]1Q[W4X2
48>PRCXb/L3;7J-^=BO(CE]00G9.+:)TV6P:S_ZXM6GS^#(G+D_ECQD,Xb/;P^CN
gWBD^cb+2U/b,XL4YDAQ66_VV/XZa,SD)^4E<,6D-bL#Y+XE[.W2.9/eLGIENFaD
+_:7=71f4b1f?Xe]EJ:e.[K:f@^VJAeMEADcDU#VgE^a:Gf3^R4f_d6Bg(7d[F55
6.47^O3a#Q?bTe7U[b]YC6)LZ3@JfPb-B7Y:WRE&5gF-O_SV&GQ_9S;b-.BR@3#S
6JZ\KVBcKY/K5Q2M^U3,\.e/A[^a/Jc8[<,>[<PZ2[Hdc4DH7@+#9@)H8TYcPJe[
N[e)Y<eXXXB3.MEPfE2ARQ+)M9/<O6@DR@FKO&M\K6G0@VAEXK1fJ,b4AXM,(G_^
?.62@E4J,T;^-9Eg:O[L]&Y1gc72#[a,F=2K&GT4KZNSR;dW?B1d(9MT(=8_/)U[
075MY#E^Vg?gG0P8]P[.OM67DS@I2<>VePN/W[)EE1/561DNbI/)U[M;V:d.IcK@
>C>/Z3HM<=9MWRI0.D,P6GcWP<5E95\NQDZJ-GcDKP-E/L&[=eCF[[&@cT/G@RHf
+5+:LcXYMTbeG<7@30K?+IRe=,3Ab,L+])DIc1GaMD,bZY<4O&_O\<=O7HH.;;EM
dIb/@O+_<?RF,/C:(7f[BK[YZ16X=>RX=T&-B=UeVGUC\P45M:N#T9V#DO4^B;XP
/+0,5DWOW7>Zg?V8Wc-AQ).U&=AaFRS_W7SCO3KRe&,=DH/Xd7WdN#f6JAZV(fS^
DN/K]V.[#,>dN.<,NW)]4^6f<fBNW]66.[K1][1TFd_&0Pb2Z]d]?I6TP(Y,YV.c
5FU0S&QHX?-Qb,d8a7/:].;<Q6CY:D^PR+:C2>D1ZMPSV2=II4@.3bg2)+GF<4[X
A)(dH5-?3XV1=KKB33G0:322H[,[C5\g368bH]P.\Y:4HV.e_((^[UY+Ngf6gT/7
5N7(E]77Qg=L^[2Vg\>#KPg@2GG3FcgK2_&<UDFI1:XG&]=90AT#I0WA?@P#62[E
([3PRX,;KS?b?#W35ZZ-K3NXEc2)&=>S?.0OQG3a_ge+B80DXd_5,/>X=:YZ))FY
LH8_R.9d0,>\_<L_Y#[<NV0<4=<?Mg0X)LN<P[CL-L2X:EBP9UYJaEE]Q?,PWPK;
I]KO08b06JKb,,X/@M\fUS9YFcF294>E,BAS3a,1(937V[V,18=6JY=\34@d)XN_
0b/aX\\##_20[7VG8X9>VHFN:Yb].Y;R>AA,F@N.cb059eWLg>9dYa1/aR?#])BT
MN>GaAM80LJPTSWaRSF@\AU^D,OAf=QL@Z:#X)2>M2N^8AW\ZIS@&<OC/feKUd2+
1KD_\Z?6&L3[Q2E#U\<A5SZTUDR?78QI6\-74&-E0Y]8L@_/S+3AS=.#]gUG8C09
3UBL0e+\;4R^;bAY&K;4C3V/O?Zf+>CNV3c1I&)W3NWJ?DN]6(WCOK(SPMeWU]/4
WUa-F<XV@[VXI,fE4e;7R<V1_I8QDX4HG\/U2C2+C1Od/Y7d]:\N=Y&^9/0GA6Oe
,-KH^0XW(UKA9N4X.TR)L5C.(<?-.9(Z;5e59U><EC51LB(H0fa9E-g;.SH5IO8O
UL57&^??T>VdFZVg3>PCMQc9f:N65Y3-dQV7=];S;]EW)/a=9(W5+B+[bLEG3Df5
1C/<IGB=,6XI_DaP4#b\2F0ELFAfY?3?bOG;C(I?GMc=D&V]D.cUTA?\+9Gc&Gec
AMS7MKI[)b\LCWQ-KP:2S2P^T(+1HF[3e0((?-8LVbbbQc?_NZY=C9R-NefC8[(W
=-B>B@De/-H678a2?68MC#3MW)0Bd+H#a^c31I+K4b@a+G,gQ?dW[>P^19,Ib#]^
Va57EO:>>6_Ec5c0d/6K&+>INDKBd0]CabIHQS<B=(<?FJYQ.+<8gVQH@7WV[]0(
3FJ3BQDZN.OK@b#+RA-001/9KJ&^?M+G^KG4Yg]753IT4)BPU[_N3fD\0Igc&@PE
^HD5[?]GYTTDMO.]<<fL4_82TG;GAH(L<a5bIRIP>S@:BG0W:X4da^Cg?YR&;)Xa
1HSbdBae/1T9TH<d:d.#MfHD7K:=<H4>Y23I)>(BfDE56W5)D/-[-#Q_0#YJD<c@
\/=4D)VUP[(>/Ma-?C^gKLO-?6f;a3S._=]-Nd93ZIC9Xb\Q#^:Pc(U2T>96_]#=
ZV6-dAd,Q2?U]GgcC=6[1(]@_40BV)(Pf2Pa(GAgC-#;3>D\f.Y:ORJ7TO70]cVD
>3E9V=T1N4]?f.FFN+9<I11=\RC\0.\Q2UXUO]0^T>.UX56aNA00;/cIQbECZAdU
#daZ2=A<U8B_O/&SZ-28GDAJ/<gD/VZD=dcZ9S27P.M6@_(Y-Db4@5cTgD,U4>b(
Y80W4PZ#4=dZD/a:F8;;=87fRe8460:S?Neg\GJQ<F9=Rf5:33<bHL&#UdB+?gJK
BQ03\B/QY^5H+0@Ff:V4?&cTA,NP6L\MUBQf=[;Nc=4>60V&X_Q_4Y[6)W^bZWMa
Y&JYg6F0Y^c[d7,e@.bHEM5JN/BZNE-JW+^a>:_NH56ETTL[#PH9^Ieg0<gA_FZ8
J-?3d4RX3\e+c>H?41K5>=1g,NL=6P.C;+<d]Q+0<#5,<<KOYS=H>e\B1AK^NSg;
T^2)/+NH?aY;UD5faQaD^1W\_2(N#5c2,=]@-O)-DV:7f>[XG14A2799U?<EeM.#
27_.2X=\I3<<Y,HI\2E633I7I#/HZC(JC\]?IZ/D5V>7^N-L85@f20^7bT6NFF?G
<CdS<,HJSP?;:c8K;.Ecb-fW439610F&YJSK=18D8#8;/RX&#.2S=fA5Y_[NCSOY
U++CIT749+3KHfCLJgX,59)U#TQ2[\80J41>]+H4U2<=O_(K07I?WgM8Sb@?SX)#
.S;UOP-3_FE;8f-)\O=CgINZ]-Za1N17U+A#bTFH&+.)5=[M2/+KEIMb?aH0UTIG
a6b&XWEV:_RIS9B;CMMK==78Ee8260FX(b[2VcJBBO>N,0.>+XU;UW5Xd/@[MD<1
@2S50D=d-(0>d?&^7.BGCe9?4K>Z<2O&AUgAI1>5(Q9^JRZ4X5@M&,NVSdK&0B[J
N=5[SZ.G4=3XN122(Ld#QcOKGd3X(_T7Rd5JC)F7Vg+,+2b))2EJ=b1ODUGZF[5-
BY\UD48e/+/Q;ZZd_D:C2O.6b6[&<NTM;b7BW/ec4T-,[XZgGECBe0(@YNB=PE(G
8a<e55c#7[?dM+=D7(@/Q,2H<9b;Q\IIHER;FP,&)_UW:d[+Y[[,J#N7L/=cC+e]
CbGMaD>f7UWGT,>QAIR9b@f_^/M46AD:8NP&\1ZBJe(?gF.:=2De#WBKMHP/-C/^
B9#NTJW2[NIH++@Ig@/;)SQd8F_O?b^D8P?C8@7\&A2.5D:gE3N+[@gZYGN1Z;JQ
#:I992A;_DY]B;1W>_W?)XH1F/aC7A&0-G.5S/QaXA0>E)f<5_W/K-P]E=_f9IHS
eXA8<eE3\D4Q1,;K48Ee_MOb&]6<[JeV,2\H)1#EOX1\TX<1-:M#ZS4FIAMP#UOb
^S,U>CV?VaF=Hc4N/,gUTQKbPT;8]+QIJ2N@F4dH-;Q;E=Q2]aS/[ZF?N)H\Je,Q
Cac[ND(eLC/-_fQa)d;gcBea>gc9BeWH@/DHA/#a]6O/aKe0.EI:#_-8d_>f89(Z
KGg0P(0DUI(3.DF?a/eDfG_=)MHZSEL@a,0e4CLP6)&KH+aD.f1^NK-AZ8KIa]M7
M,[QPF<UYCZ&R&G;(7@&8Q7HgNgf>FR&Q/:=MLS[EBE4<]@9;1M>ET:,U#=.(?:&
g#)]+)4:KD4_R[0Ja<QWbba8(4Y/P_ccBHB_XVR=L.<F<-:?T8Y33,:Jb&c@b\@8
1\fF5UI(J0g?2[VW69A=gJ-5N1&VP][fc\;2E<:(YUV3a:a@S5@g25VRG6b1LeeX
DD:07))^1,]3YNgSF(a?<0cZeS\1bY-#1X<436L.R.70084J094X417:2UKRPM=2
]TPGeGJ3f&YabTcB\@1K@VJKc]M4-C9d9^\40X0CNZ>_BTEeQ+W&J(X.ce^MO/&Q
a2<8UdQa.R2V);X5@YY]#H-F0(,V9JN2\IA42bVHc.\)9&NVO?f#<OX.@>#XFAG-
BPY77+[G4O9HXR4OXZ/?PSH0+I?T>^8@>-Q\F@XQ>\U4<)8EG5^>_W):JWD)/&_f
3_U]&T(1[R6#[^D3HDc=E>T:9APKJ/<Y4NQb6f5@R2E>Q@6f]U+;)212.&LAf/bf
YOPL;\C#NYZAcU4_<L+UY1:?MN3\<O.W\2eZbWO9S7HF+]+g9c?K49(Qce:CG8];
4<H4TA-cWC^c>:V(W\VVIP8(OL2?fg/c7\CWI7&_0/2fTf^]Ef^T9KDLL;+S;RFG
H#ZfFH<Hc/KQ,8GJSTR;FEO7L>6EXVN;Zf\7gJZD8^0>SbQTA[@a@0;3;7Jb,>>#
\YG/ZWR1DOe5EXP)CE:3XD,XTCG&9Q59R4^>VV]G?YYSG1/TBd@ZX\V=OT\5-c1T
+TWcXL<Y0L)b+b5ZD@;B:UTWK_?3[8@F;ZK+Z4^:aM.+>,&02H9_V&eWKg)B\dA0
a-\[=:IH?:WT]Af1Z)H/.Q;QU4C.gW=9P5+g75Yg7d^+Ja^b,>D8-&LP0Vb,dX3/
Pc0NW_&QQ2.#GBMJe)6U/](g1;L0]S6SQ=W=^V;S_5_\I1bf@4N#=#=L8RY_d2cg
OeGQ&Sb9P]UD^3-[gQZ[^1PA(\1R#X/<BM>;8X>#MD:&P0PJJK/D[^.,gB^f_O?7
F6^-#9c7KT+6LZ&,c:UPd@\Cc?E^AaV+V((6/LNL_B8,c4..FILE&S2V[f?R45?G
6D3C(ND/WDR9C5[3&G5.8]T7Qc(FUL&676T_6=WJ[PQBFC0CE3M<0T@J]c@Cg</X
)UcBGUaOH)?F^P1f?JZ<2,D/bbe:XVQ^OTBC/S,[fPX[8<(N+BFTV=cff>D#N-X8
J\30NX4Ra^3b.NI.4HSP?2Y<FB<\N];JIG?S&>CQ\6EWC]&+G@>MV/+JT)\_PMQY
@?>6MI(98>TOJcXU:Ra=g=ZEEfS<6#NTT>ESd#C8(DR)1&Wa-.Q,&fYO.>R&c87e
MbT.P3cR65D8UMg+FbS;#:CG)+6Fa720>#XLWOf/C#]MB^ZeH@3(dD?CPQL.76A#
3(Md]@N+B<UDda-&:E.,8COQ@XOG^]D6a);K(?;Y@GP5UG18M]6(3Mb5&2J0c.IJ
@>+SZc#H8YQMJ;E.E11.AMF&K_#>Z7=UfE-PY==a7.a#(H-Q_,752_D=;e7dQaRE
A(/a?+/\)#528LPUZ?ZLa6G6853S<gDg&0#LU_-_-]A&&[U1=_/VW>\HHMe]L6-N
GT4<.^a[bDJ2c0EL-E+42O?<0aV.T]QTa_dJ\Y:JTa,_YfB:YEfcM1-4_X)R3HG_
6;\@e:acX^RSD;2GI:fWMePeH=bD.6D7d1]0GL_>P]?^L:cJ0:E+2\0<+;:YWHcO
MJ8FXQEeIYEM?cYF(Q6U7=Y#9)=)aMdB-B@eM+I)MF?]ZM/ATPBES,MH4ZMD)43d
F8D@HQS6d2b)3_RR3HKa7ZLfeFe/6I1\)HWAg2=cWKS12^?80+T7)d:+EcE9gW2<
]&J/.Z#3Y;DAc;AMVJFa_&-3>@,Ja#,5NPN^036Q+Q4A>Eg@<HHQ:UN5b2LDN1@1
B9_L[)69D5Y#?LX\MPXa;S?R9.716X87(VX2:&<XY4U=g[>KWLDB&IP?93f,[8Xb
[P&72Cdc-d/_6,8cUO2)JefNM]@TT)3Ycg-=/RAOfQTDN,Q^8;g6Cb<YB4]Q\_/F
8U5e(QL;41?V;CK]3aA@U/OeQ\\<b8]S1e88R)bS@e5CA@IH,P)+3O-YI0YLI7,S
UWE,E\eIM4O2M^0Oa#VE:OG2;DG.JD/W;Eaf,S6\ZMT?TCK3=?^_Of]V&6U]SGA>
X;9Q-/15TH-BMM9g+XP:)+EH?3JQQVA1d-@/_HPcTgcM<H79MC.VE;A9->@W60DZ
4TEO]J.,U5(BW8c#L&?BDAQ+#^gCc?0&0)Vd9(#&\G>HJ3QQJ8N5F.N1NaKBUF1@
QZXd,N)BC;@ScH/Q7+#:9+-4(+.(X<2V-CKCBQ7If(S8WTT=13Q1e0A&\VBL#8=W
GD.0\LMeVc,a<]8PeZ&QR:=2(DCfH8fSFIRT&9/XL+>^@/J9/ZT9XKU;/fN8-+Jb
R&(S1Q\5V&I#_F8;;=fD^D22gI^:OP0CK8WNI_LVK2W:FB#7-6Z69_N\gFDPT-IY
H&@RC=2Y#RaK:8S)gVUY?-+79?a[FgZA_V[BM]2PD:YeV1AbX_6V0FCS)\P)V^7>
&&^40G)E8]5&GU[<.[dYMBXBTKS6aR@Ve<=ZLaWS1?7QfL)YM[CI\d=IbNbeU)#\
MB1PHP@DO8L^D>^>B<Y5_-JO3AC]V25/a,#I4.,2c6OL2UXOK.<UQ1LgJTD2:]99
CN[?b7P?LJ=\OJBHJ/+LM1CC?;=CaNR,W->A[1b<1<8RR[^D1(O[JQE5H\cb<=N2
IKf0=:<9HL@XffT+V<PPIcST[BW.=NcV:(gUAd#gBO-G(fM@)+[3>Y-+DQ61OX4I
E5;agW><L-LH4M=#6b<4eR3^]\?<9_):]fRF55=^/4KBGL_6]T1de)[K]OV9HQ/D
J&;2]EC3Vdf?LI7]5CVTbCF@X+9Ig-OG+U9U,P(<TW1f>(VF15;.5-O29H3P?JV>
Z==&HJK_=_.b(QG\2RYVWX=:W21EfIg4.bAV?JUgC32F/,OMO_GO/:DUaXAd3PM[
6LNZK9L6M(9WcDS.P8_DN1@1CD_e:^K3:J&^C3SMEa-4?ELYXV=ZgO>QS;,3/+;C
L<G=,?CR[cC<R1gJAD:Z9&=)4SXcP7QN7R3f8D#f-dITSQ9VO.D+PeH9]?6g>d.A
5Z7>\]VDV9]fQON^]&#K?G0J)43<@9&97Kg0Ld6geD]W.QfJaH(dU[L?OJNT>THV
cGVN?e+/.Ic9-=[<ePB?bU#NA)E3L5&F9<#_L1)L^0>C8I2C]M??&?4GR8aJ5N\,
g.]3TG77FOUM)EQVSA\1X-WU]2UNNfX^b2WEN[c3W_a@c-N0L86;fM&R6[M[UYN,
.J3(=@,e)[g&#@Q(dL/Q>0_8Zaf7#P((=#B+,G)aA2#(3/&c4NMQMdL7HVOHcfV#
2+Q;_M9\O@)Y6C@5[[OCX\NKG?=\RTOM<BIab[3AgNX6[[+-31Q:ABMcJT.)TIbB
].C5_RP(V=b:OQ/KC7?9J(fAN]-9G0bR&2/I3?(2JX.3L^OV+1Hd1T+#QB_H\V#N
]aIR_I]S<)b\<O7WNRK9/a:/44ISJ5Xc:HFYLA205#Fc<O>CP,(?BQTbXd(a)39L
,?)I:6MIa,CDB5S,<(]VT^OJ1<<VK\BZdVCdI)0DJNQ(gXf9d5C@b<E<LF3Qb_E#
.fb(+<EfPeDI>bM\G@RANeIMZ[g9XFZS#RfG&,L9[#\\FFVX6\7YXOE-U1;64(cH
@CaJd9F_+&02[><?RYWS7U3(-=4Y>0-7cRC1YSfTUN]3B,CfH7M)W^IK6ZVY>TTd
TebNEM>>33W#cSQ_.N>_8^LUHU:1M7#HB_<?ea;&XH;4NGf=G)P6<EAUb683.RQ-
WKW)3YK8@[c.RdN?@74gSJ8B0<BJSIHYeMT2ZS\-[4RcbO_83(<9,d3])5/EXaQX
e<C(X)W+=8QL@a/c,>;<8D2cG0)PW03K[:&.BaSc5\DNbfYG71O]<=6B0TCA>[BC
G\>SUAdHT7/PQ-+gaA/WeBNbFEFQ+4P_(SZaaFfFIb+f4Q5OW#ceRP9+82I2-L<6
d=d);FG^FgD3.X5&Qe&I]AH8KSD)<<1I/eKf9@7PB>/,NL)B7a]MOTL0=]_7-@#e
D;:C=KSaU@O9Q4;U6gV?ZROFB>g1B8&gg=3G1H?T>+#c4H5N=E70<=49/\VR8PI:
DUL6O_7^L.Y;S/IW9#a\#)f,[^Rcd36GIM<0N./=S.8,0@aBf#1IFb697,=-5#0-
(.3Ca@cH2g/[A<7cbgIO)2R+L?5LZWJJ.]d?I+H>U8](1U^SL?1b\/FV2/a9E.0Y
\I+I.<Sb,P3\SCFJfK^7^?UMOXgbB+F[G_ZG66\Sa@BZ&D.cO[Y,^]AV.ScEZWNO
W,bEggR6MZ6dZ(g;5_]<;G1G_F9GcK]D0TJPEI@>W)?9NOg]3F\0O_6aJ>RM[25E
Y)M_Q8].>aJ-CLQcCe=ZTgb_CR6ET8.?Q;L^JQED_3<9&(]f^#59(C8V<(e0?=aX
9g1\X#MVY<=J+.fc-P]@^8\7J_cYQbb+K/UQ\YX?R1>\,-&0\M=E3)-R1(&_A6#U
I>LFI?]\?K_,eA4Gd3@&DcJRSbfP&\?/D7OB-6:V1#SW@Rf7Q>(1XB/5FWdLG88T
\IQ[=&dM<U74PZ^.<W=QZNIT<FI>eU@60))PFNbNO6FPgGbG^NGf/4NGPc&]XA+f
JDYW^Ig3+.0T8c02]cXVH>7KLZ8+F=@KQPM/a88W4Mb=JfCW^a;G,SH0][Me2KZX
KUeH4?0IfY^P4E,WffH)T[90=2^R&E;B>66aM.6ZE[(A)=9LZbSN>>Ob9g(-252V
f/eMB:TdaTF)IF-eJ+BQ^4:=5Cd<V<&C]_GS1R7?C2A?6Sb\Z/M;P[)MIO[2S2)X
]-U[eS<;@0S;7S9+WaF1,3>EJ^?R0.-N<?SFb4KC/5Q=6I],;TZBDT\[+b0)WCa>
d60<A;#eW_SQa(,Q#7P&@>-C-f#Z0WP/#SIe61MW,fd_P.&^3LGZ6>V7-NR_)M.&
G2O[?J:-Yc#^BWaR5:-W]Z-YWKDL#VOCHa#aU\6=^5<D.7cJZT52Hg8#Oc91TQd;
ab9#G=7T>I;Z/LYQT>2VA;U0#>M\B6@K9=&)@c<T99YVP2]c#6SGH5FP;KaKJ4-_
DJYdL0XNZUSOLZGLD:HZB2)[UaS-)SGPQ(W1KUE3G>a>4VSH,\+a@P#?V;K(M6PH
2&#gX0E]3925>aBN-af0@G27BUT-X/VS3IB)<JM>Ua^\V9X2U014f+e=fUOZ@bX+
EXM#ST)Z;JWB>-\;L-(D,\4B(N9+L?./=X;;4Gb_BF3;2_STOIAa\((W+&.-@IKS
9PLE@DBZ9#Q+>C+V=Yd4+cP+f@gZ.XMbN49)g/B&=GEK&cdBR]4QT_VbWLPF6^XJ
GaM&G0[-@a;Ue^]8903Q;N?;+I:01_;Ea1NbL&(bZ(/X(>?KF#ST/7^-F5K^3M8d
8.gH-S(]=BOX0=PJIV;WH2T_[G4I&DD9LC]a[-?@BJGbG.R^TGKA]Vg.6:Y+;JT2
RCCC1VHV@EQR)#[X.-^gObe>XN7H8_M<V=eLO7D:JDVb1L\^16D/D@(&eWeNO03(
I6V]2F9C4T3=f>EP-?/T2Lg1/3c/:H;_Q5dE;.^3R@7cQK8&[([2.NK=e=(VT]RI
)\WGK-2L,844@=,_.@]=b:VB):X6UW6.NMPVQXA<\\?SF9-VT<ORScAbVW((^<gf
SBSIf]c3C&0)b/DJX4)TU;g3^[ObFf3>MW1cZK\:YG3[D19.Q&DaTe__/@gc4).P
A-I/K>;K:\[:2H=fBBA>A=Ybf]J,4S(gQ9J&Y0Ff+D>O.;B/39\GFBcda>2-d38F
1L@Y<^>FH>D5&Pf4g0d]JDQU+(55=QTFJK=&=99S=Gd3+R&a-CcgD&C\W<JTcP7=
YUY#K.1A#GR(_4@.+f92>=CJ3fa3J3:GfB^=D67R?1E>B/^b?>8RZ<3(K#=//^:J
Z,(L#IO6[QC(NY:\-(#3a&.<YIA<H.J+?B<UgCf\WT)f9?Q(W+X;D;f-eG,Fa\=^
VP&=cQ7S/ce>dc>RMa]5L(S^_./.DfHAH^NI3S[DRP;-2:YgeTH>CbYXd5)f2E8W
P]DVfGKR62bSF>[ZOd.@^:?TH_1U&=@7^&-2d,bSRJJRg_@V:R3HB/[Xc&P>aHbK
W,,;NfcA21C>]c1MR1,e@5XE^)@=L=?P9T<3SE>DceaNX\9?D?^AF7<>Fa/&AGSY
/^-C8AQ2,BV<5c(4]Vb8SC(9TEX;5^4^&<9S7LH_L#eMK_AF5UbLH(e;AV=aAU_W
Q4?H-/=X\CJ)+0T/:1_5R4CR+f)Z#?AA_?TPLC/W<)XVB_US7D-++NMVGNcU^eSM
25AZ[1OgDNX5;3@A.1I2KL?KPOc\3T];#eRAV+SND>fOXY]0/1Rf#RLJUC82DBJg
S]9,/1[+Sg^XBBTFZ[_EeBc43SJ<:O<IZ:5Y6MG/VgX;[^Z&Ed\FB/7QX\#FV+,E
K-7B81@;Wa1BeSWI&09ZQ^^7E;C6Lb=N&&dUP2J[ZdAZ5[O:bYdNA.,eZ57#BF-6
DK\\H[;U7D<\S?fB2>HgdSY_DA1X4L4GBSd=0bHQA/=L8[U)HXN)FcE^372V+-9\
#eZ)-KE-X)@>+c:OQTUE<[F6+0(YAc\Z/MG)V\fXc.?=6EDR(<3)Ee91(2;NCc@G
TC9aXY)94<8]-c);bKP@>FEeD</.CC24&.DCV6CD8/(Q:PgW4,FCV+ReCS[).)dU
+F^XC\7&0N.+O.+6MHM3@3C-/BHD)0OS2:XccPF)^VO.;3-(/B?gWY7Lc)/aHC4&
Z8fU[NAZ71;_,W+7F&<D#9>Y3+G(P_P&-ePb(-U]Z,[8;Nb06f-WN@<dee>K5e3g
fd7B/1?KQSV<AAdDG,e#;<HX\f9_b/-CMR4YUO7;3#29MH?MD<@X]c(;X+]W=S[,
@=AAF8A314:)a]TCcFLPP5<)T6#ZW_7R(HYHQ]#NaCPAI+KG_Ee])Z&2>OFO&5>X
.d0=7;94)UQ-1PF+GabV0\X9PAH_@BaM\eIdc^Z]Y\X?-2,;c/Y?cHU;b,BW3d,R
5aNF0H+Vc^96-R3Vfb6E?d42.bESZ5OEL/<+J84Rd<;\F7N^-70BGc.f0W>(=Y7Z
<8B>>&.3U+8B>L:aZ1BK;YaD)14NfYb8<,Scd[E^f,-]7>cARV4(OKXW+-D:57D#
^4cNUAHL@XC?0f>?@aF=:WXf=?50/IR#9<GFdASOBUF1>21VD?1b(-fH+]\[a?FR
/Q>DM<([ege>9^dFTB)2]?X=P4)X7BE+^1PTEf;fIYRK1Y-&&:A#1VW>JfH-D0NF
^c]7eWQ;]KFb^:=\X]c:LT-J<((HAOf8b?F&IOB.F:EBPBPSJHS,e>[[S?5:GK0)
e94=7@a/+#dE]0Y&<1IM?g(N,\7U.c@\/BMaFY9N>0A.cC?N5W=J[8GVSe>\/5Qf
@6^5#V_W2[^#LYO9P:_fX:B3VXN)NAa5ZfO=<M7DP-A]A48F@e\7N/3cG@O@,O82
LacA_FRW3P)NdDBcA^IMg/Wg0bdTb;S./B-(M+aUOda6bb:5Q:(_f\-;>W8GQ82?
gc@O&)+H++^R)DUe_/#F1SDagd^:5RQ_Ac8?/N+fM_Kf4&CAdN(?@/,;5>1;6c,7
SB#AD#bB(+GSP_Q_6=72]E:Qa2WNC@2NY6S;JdG(^(FNYTP3IUU_RHQ,E>cQ6WE>
5CT6_NYHE6-;?XEbG.[3GJ/8(,E5?[_c>B8eO#JG9)g;).F78//J/</Y9c)##C+J
72/VIL]H28fG5?H_1P[CN]fZG@XKa@e^/@L:d8+e+YdZB6N94AGD_Z4e8^_8,?GU
+BB(eK2:(dgBF-^P0Z#,W@Ka-LPLgS@FGKd.FQZf<)KLIdU0@:S=FQ(&Z@P/d+<1
;Kf/D_519NYW(#Z1aJC&a7=^4cSCdQE@]@,J4107A:=6EC10Y6?P&Q3BRdQV,Z4=
Ke5EaWVW>D>K.IcQ+R6c^]Y2#5VH^@]+K7-f:]E-#?]U/P[VMQ;=/#&TeT[fKK[;
G;>bg?M.Gd>BQIaQ+Sa[R,CR[;.=M#&f8Sf(Q8V,(<TP[W3,)JG/bb/CY2N9Kcf0
dUb8Ug?YK/;K+M9<M7.d]M3SP:&_N(RJ/BMVFbO)UZE2166O.5M1L,^)<SAAXd=P
\:RZE9N:TF8aVHGD7f6#4(fPQ(<N[fEE.\8:)0P0/X(@<7ZI/(H26.19_W.caU=K
E[aa#&/6NCSM<WA[^E]1\^)Me7V-S@ZU#KO9GPS#5:RL<Q0I8LL.<Ne<#;Mb0Q:+
_L1G>OY]TJW,_>PC2[W?DT&[+a7CT6W4Z_TZYVBYUd2Y7A\fV;b1O1[0NOOX<?/_
g@HUD-Da0?_QX&MJ:-GJ]EE;FVM2/aZ\c1;+]Tbb65]QJTd8?VPI;d?\dgCZ2c.U
_CS#6YTffH@<4O534FIFfa?^=e:PfdOA#>Y<S@65,(2M0V<B>AK-7O8AfO?Tf)>0
\J&W>VJD-,K,^=/EdYEa88AaCDCKLT<4:aH:Ud8I)Z-&C4X8C8+VR1>:MB6@I2]8
e?c7:dHZTR0ZF6eA(QfX(:7<Oa2+[S+7bg]<N?#:U_HRY6R7=\;KYXaPU+1gWTCf
DBM4?.Uc]H)3>)]7<\^H0KMO4-JP2YRA=SW;UIM@?X6041d?4DGfRDadQ)LR0d=_
/1XZe4_@^ZN1V09dKbe(MSa/f10JJB,F#JGO\L,W,Z=RO<F,V(Q\_6DK,?(]AU_2
gTQE0KQCAA34XVE)F;A^-#G\YfcCRd:6^O./-W(D]1MON<P,Z?d@gaZI@:OE2\O3
?&/T[NKAR)K:/OG.DI&8ce0^-X=FQbMEf<dB<?:a:9MZeBQcR5+.b5=1e:e+<:&=
8V]\7ZM@3:L?cPJ&#>T5aI:C)9?;=]OGL(Le,UJf11[]^-]A6&/Y6AM;CAadA,36
K)V=.,)I^(C76(Kd4GH4P&H)?6@1X=NcS&-bOQ(KA]SU21JZAMCGa]R];,BR8fXQ
Q]AK]^f;?P=KZ)NA<56[(#beK2f\0&3C0B>S5c3@+^[(^b#,KIVD=\Y4)4dQ5PMM
+>GM?DD[g(\WWQeU0e7.S\_48b)L32KQU_FZ6W/-J6XFSN,>[1]a,bb1eZ;H\ERN
BU;W124KPDPRJPJ+2B_J;C3^gMf)Df_##bO=T9+gcK0NU:R)KZaHQ]4H)c/<&DD1
NTL^:P65K(QM,]g.@1EZ=.5,\C5],<RC(K0)\D;-+PJK)XS#M-#VF74?2WOe@U42
.0QbO@S++;Q][3,M5fEe-H/bB4a<Ac#?OBMI-&ZKE4C.?fD@9g&>=2BTM3E(-NWF
\\267.P6.3g([#>PTbe.X0LCAJFDI3^<d30KG>cI4C0Cg1?e[N4d&B@>/=0E&g<Q
Q6/&D5L;/;+(W4^)bRIe?C+3\/_>Z[O5A6a&TRQHcU@HbE8G=[(R)V8/R0=bT,;,
)e]X0WP7D,:JW0=LQRX2_I+:XC;1Pe)\+:0.AXWgNTCPMa-35SW:>C#QD29;;E.\
fV;d-\N1LP1UdD+CW8D,XHOGVYSVV_E8D/4cJTRYLL@/I+QG0,#R#Hc/@eBH23[R
MVJ9f>\5?UF__S]-<A>efP/AVQ^fY)_d<MVSAF7,+5UCXQY1DZIQ9_BK0_?[EWB9
Pg4&WZXBNE#K45A>?Y](O+J/2P9ef5CBb+eL>U73OO/@QO&0F\.U44LUC][Y(P1G
#f,>c_NCAE[<e[6ODJ:6<0>PaQY94E+]1_A\E1>E6;3=]c[e/[a-^:SKR-:CMF1E
C\&,g#@T;16-VEc;(\:,/ceR#cA.M=\9[;3eQ.[M[,Q6R\e,<;83[&AHE:B-<AQ1
dfEH,:RFUF_cB)>[C@](B;VX\Y?-YPM.b1TJbg:QI)UcMMR#^TV8R^6<,K:W.\\R
a+(gJ[9?OKF.EC5S43dHg5D;g>\DPcDJLg0,W3aS;R3?7:(2O8WYBfIASKgQd(WY
b[QQaK:2gdF#cCg@_HEVUXC;-^caB<8I/X7XeH6^<9@?3(R?:W^IN-RQ?F(e9>22
c[cU(68R)f29Y>D=>AP]<O9Se8;\+)+Tf-&f<>eHPLZdG^0<bgOCFV8NV)C1g]ge
DYbJWb><&,g94(U^@O^ML8.+],1[(6Z+:UC/5a?:VWWZ6]H+5\QO92\7S/Pc5\:]
.c\FUIdX=D\8f3UXB3I@^Kf_G6>3?UX9f14C4[:4_H2V7K_NBAIa0c/QQF/8,GK>
POG:M]EZ<@8&7UI(J^-J/956KbJW?5Z@M2]B#PR1J>BeL[CEJ5bBd?Fe(1#[4]7d
3/^N+3fEd3+FKLN6#4GZ-@UNGJD0#C)b-#+eSG)QR6M@#\]F1a.Z/fR2=D^G49Q&
)>UDY_Z=A?d<EN8fYQE<>fRb2W5U[YIZO<5NS5]eV@I=]>>7P>,HO1Gc1K#WTeg8
ISMGO&S\A8Pgb(f)MUC2S7\NZ6[Dd_V+SL8H^BT9FcH7XeaW;\dD-GaYRFbePIF^
P:fN-bb+SG=5D0eV&-Z4KKF8N[8^FeV\EO8.+[WWBd1P:&S4UR4;f#UIg^F9Z::B
YP&af\P-(>K=VHBQUTBCP5#)SEL+P\-V+BKeA<_YTA+2R\dc<M\ce-5QOZe9_.f@
?>[\,L^(;R+5U-^4a8H/R@_X@]39AfQAg@de?/RX^TL4VOc#Kg(#[<\_?886>IK\
@S]eYL?KHN-\(,bKcO_3:]6R5HWO\Lge)3FD7UdE=JDZ))P2KL>KI,I<JG+WKFZ3
JS,Bf]^CL;XL59NM=R-X4QJ-&8g.C]WMOeQ?[K=XRbDb2?;e9Ce--IL]=dJ>YA4_
AY(XW:HQH<O(;cW+,>c@8XF5e16E:39NBT=6-QM8UYYQC..DZY(:ZX?UaUO_Z9gZ
+5c3FQB-d(5@IJ?5)_YMXfRFO=DKEG&FRRKZa&\[X3_D,W>Id0\Cb++GNceX1@==
G6BXG7_FPEf?IJaY942V_;<5>&^&]X:\bJ#DdOR)#(3&gC,&fW4[X2V2&7]VYc;Z
?:M&Ld\/\)U+g<(@?<AKCg&AWGX#+-I;E0.HD\N&^\^e,9G?_P^b#aBXWSCX.FFY
4cWZE^TgVgdGIJHAD8SLW@Q98,LcVV+N?R?.C7,QM^IF/R;UgI0[PZF]=C4=U.H[
,6<e;>e)Wa#J)A)]Wa)10+DFg9WU6=Hcb@JQ-\c?;cNTcM6-[=S23RYD)&0cEC9W
DJN+6_bMO,b,dd&13ZYGHRMBG,\E#6:;1-#2c1]V=_6@bc-<QTNS+4]BBd;HV[M;
c:9KO[@G17^@;8LcB_&_(cWf1&CgO/<ZQ(F&7JF)f-;.M:,N.N5C20YI]dUGK^Jf
8@eXQS75OA3OAA<Y;N21]7@]e#3TVN[/]E@WNa\U#\C3eR<3AE_62E]]G,RfVgeA
^.E0?ZFF&XQ#D:&>T7]2-dNgSP#O/11d-FH>ZOgW9O7A-D+=R;:8QP>OCDC)04/B
dMd4G?Y<?EFAM1<cYG887=L@9fI,1MA2P]=J]e@0,.)NS0(S_H&X_8>ETKP.X4Y6
^<E9(_;C-;>#J?<cU19g54(V[9+W9gfZH)4QJB+>cL5ae9U7e4<J^>ST@RP?4S+C
=XBH)d.],-?/QA\f?T-7abA>KH_6AVc=>IK0[#Ta1J,/7BDZ/B1g1T\P)=f^7?X&
Z3DN^^R,VE;_QN2J-5AQN+O;YY@6^e(6g0CYaP=XUc+3TAM@+:AAV#AWE2K#3283
@G&=UE.?HAaM3(fb=T,I]fSNN;W56Ng6FR1NH\DKJaDTM242ZVXOLG=b<aeZMUK#
7:4I31e<A=RB5560d9#?T2,g1O8&0e5,ee;:B2BGZJ&/\&O3:&>P[)+J6^6gVYVQ
EaQE59ZC;)1OJAVY(gP28_Y[BKZ._8#5[F_;\=M#+^\F.c@XDN?&->f6bZYK[/_(
(RPS9G=)&Xe,e?@UXQ&L;bcYZcJD(/c+33cHEgJ/e1]QW[+QW1LWBfa+K00.QY[W
#d;Q?SZ2d2IU-NgabW<A&M6:>c]#TKeK>_9\J?4TYX<4Fa(Jba6#]<^#@BEJgN@;
4M(G@7UQ\A09KMg2>PH453@_()5&]S./P1U?QP^bN;9A4JO3TEf^/Z/eOU)?67M-
E^=FTK7X-]]f9IGTC:6gK)>7SB/OI_dNdHY8Ja9+e1@&X;>RQTW@.]Ud@+IbA/VW
>EA#(+A5cV;W7R50[W]4d1-KV>D+b]b34=3J_^@=P<T4;:XaS>E@\)1G9AE1YR9,
JSEQ5SV.Ug_P@RR3(T8c&/PGMIY?[9DPY8f#D9E/7HG;^]=:3(PEAUB8BGB^JZ4\
/,X0X7.:+/V8M:P=YG<M-e-b#8N2U\SMgG>dQ4&L;cCO.RTUH;\PfWEP.F^RaR)E
E@)WcSJfA7I(XT5_CV6gC:B53#S31,H_P[S>_Z)9V<(b>MDF,K#YR<P0Y]E?+,]5
Oe-(>S283F:VE_bc-BYWOJ\3f.\JAAY1OCb2?Cc<;.0(<[3H.^G7T,R(@KY@QGBF
=OSLJ&,2.cGE9<EDS>5Ja-cbN1#01e,2&?H@1eT505]bYWGF&Hd;Y_UARZLYXf:L
d>P\-#;)9\OTBeXKB.a+FU?eBZLe/8EdWFQFBa-O0_Ue@2E6Le]90N@1<c+PZ9F^
4S4@-,Q\gKY)T>GHR()Q]8)D=D2XQZL>1@+U6AB/LFXZ,D\]XLA50/2WK3OcTEJK
1U0V09e0>[:/ZK9#\?ZL#F/A=^<SVD+gH.AaX5EAV4)PQ1c)[M_/PTD0fWE4c0\^
_Ca;U.&Y]O9XYN?;IFGG>^NFgb1d&:VPE;[YL4@HO7+bZB<\ODE@.CSf<R1Pgb_D
b4-UO+M>,GXQY=3D1U003;>TQ-&LS^]YZaX-5-K(_=DML6#D[bGU,8Sc#5-#(/f8
#TMQ866c&]M(^;^(R1,SA3\1.4>CU,O:bIRGA8DP_J?d8M\=ABfg6)6.R,JNX1;.
U+LIS6FJC_OG>55aA48T#);]KC#V&G41SG9^[@dCa#?:,?LPb.-?I@[N9NE3:YDG
ZJ?>aTC->ADc=g+W6SA,W(CNRL3bH52R0&/(=KK,.YUf61.Q\9GXOOQ3-9F@2FUF
_YH8/<7/aV=BR^C3V3VBgA84W0BNF?J4CH=FIE3D_3H3SVEZF7I:Dg9A=\W49R3c
6.XSFRLE5gbA14-+f<Y\YP)fX,IC3=35Hg/ROKXK+B::&DWd_C8+3FEZ^a2R&YE]
)._:3)KBbWJ(TQZ^YCKA-bgPcJ:CCSFK>5#4KJ+0RM3S/D-0Q?)T5=GK-3,B>1V3
d8?B6CCE#;M0Y;>a.3W?0FZ6\,Cf1L^e\DI((9\_/g_S,>M3[^2FOQC7J4d,LQI6
MQIG[MeMKccT3ICV)L?-C+C83Z@GKccXTVe=PI&4eNS122Q\?[TM7MdP2:VCJg<G
#Y0?a;d.d):-IJ4^1E.5QKZ/-&:B\I>/AROc[_aD>0_PC2I/E^];.MT;8F0WK.-f
KcZUIa&7PdVO?c^G3f,5_8FcZDU@Nf+FQU&>(#U10G1_3&SN.I;J?@X=2)_dM)I.
+g@L7?5EM?#aA,/d>/<5;7#d[R1X9UcS;S/F^C/S3U@J8PeF@C?FQ]faJ(e-M^77
4W=Mac,YS)^FR]#29b8N)]<[>_.JZ+-X>cO.d#IK,.g==L_US4O^Y18-PE:?O_g9
Y0\cOg;\;2#W-b;DfePKZeXbDK;e=/bKHEd^PL&2&fQN0;8V(.DFfHMOf\6SE#\@
,<bEQf^L7+C7/3Z1ffDQ4)0M^=ZeCN4RFf6U//aD3]:M2?(B-Fad5QG(A@VS5DH^
C.EL:60H>C&\-XWb>FDEC<I/2XBV_(<)K)d+8AM[Af>@[]B]_ccK;&NP4F_)JZWC
.[U@\[;2.a\)6eW,[PI7SMR5[ZNFIaGcAFcAC[#,CB0>QS\+<bSe],:X@TYXIJ5P
04\UBDVL+6N=GE.]9FKfA0@W]_DI\]UK)8,^V+eA_\U++GMZCdWQfB#\aIc#JGLf
b/)1Z..WXJR0RNMA_fFF8=LYQJ)[OUa07G4b,MG3>#g2=Lc[_a[A5)W2Z3](=CN>
M.CL?ZZ;?:g>bJ5?8+B]=+73?SD4<7fV:d5/16Fc\U8b]I^f]0dUE)ea5HBTgYVU
1CSD3I;.d<AZIDIQR.SWU\A3\bHeeIM4=gI:PZc(SbBZA(59KSO<ZC/Bg1Z&X&=B
7(-(:AXQfFb?H.f@&\]G06#57+-@bCcQKKAWMWZR77:-U#ATMI-FTES?d?8KFgH.
VX,X,Q/0?>@_VV2bL<+[AXNT0Da<NFB-K?+/B29a,BBd1eJ^a.YeH.082+.-_N/d
fC1;R.Jg]UZSH=?0S&MJ8bRIO(_W;Eb;UJEf7&)Ta;4G=S]._5Ac&<J4<L5T[4M(
KUQ1Y#f46cD,IbOgB#2#)D)&(D5;9LY@NcZ][fFWXKJbP/#gEIO);g0KDT^;Z/KH
5P7/PW.g[LWDDK[C\W51V]0PW+:/CWg#Kd8:)Q5+(SNDC[H<=PSLMgTc+EMFc7N?
.-V&WP>ULL-XV03T^G4JaNM=PF@#5S-P]K3Ga#QT-<4RAQ_&Zf)IaOTO31I3E12b
A&0B\b2>\(?B2^CWC1<X8VMV0:_+Z[bMSaROJ_.CJ(3W-O?/DgV/C[X9bDbW44ee
),^+5JC/Hc028).+7aX:M#9==K8[4LUN&OfQDL0[IA_+cE<2d4.EC8ASB28\.)+F
EbO+QWVJ>4a=XQF?UR^BQB#2=)KfM]11YOVKV01#23;2LR)e-J;:0^T/dNLQDC<Y
MM9:_/T4=?MDS6V;UCI794&O8=0?<V=U^70<XNQ[d.N>;W\1W<>1@d;WMggI^0[2
,Z\4+QP_b_)<cR:7A?9VJcG5&Hd&KSRVO&XXKLV)2:];A-XKGfU2L2N9II,OI4E8
5@LC-a(-3X<L<YT9:2E&>efMQC2I>;\S>B6+OaETd>]M;7>;]V\d_8^3a;<,[W9K
Z9R,8DWV@US<41;BSGgf/ST<VPgAVNJFCB45WbDHFKfaf1^WCM?1BG:dO8VK/f4<
-.4^9UAJdWIGbR]5K#Z6dY.WH?X3\.,2T3#_HARK_OeX,HW@^950LW2FVXZNSTDN
8_ZA^/^&X2H91/^U8X(Y>7/6G=P:#8RNP(LTO[Q8I\N7;>5G=19GB@e0^&1IF:,2
0gY7>AB89Vg1b/G)0_U^.OPeOV?FV]WdPZQfU3PR@]I6]7MJQ<<d9V^F:C]+1MM@
0-K&0#f;f<\KdK(DC??b>;B0ERLL3@P-IL^(PL#;T<)Pd3I?TTd6LT5ae32Zf6?8
Z<@b&@F+BO0)\6Kd\N\BJbRWe7V#Nc4#fDQ._g-K>YWON2888Me,S)<fC7B\LYHM
=_2/G;?\UF(>_FX45B/ea0;G6FA?/#)3b8\0&eW3^<RR+V-WceL=cKA<IM=C>3Ne
^:e_Xd&8NRU[1c5?g;46T&JTfJTKZ702?K=^U)3U<<f97NEV^?_RMOCV0HH6bIV=
SNY-SWN&UYXcA#+J0^;0GSE<1V54]FgRT72^\Fa>]KfF02&RX8##^OX\8S.0)<9;
CMV\[T(@>=aMff<B75MKD@Ybc\[fQD<L,]2Z02c:6d<G<ZL/UYV;.c#,)f2(eF&P
b96ZT;PgI7d]8+\6-I18K(Sd-)F[@JbXA2O-gD;UZ]X\H@_dJOPfC\A-4D4MSZ]1
D]/\^.KZ.V.#IDW1<?@=RP5,^(,dSKZVTN;0&g5(3Ea>1_VJM_O#L?0Nf)&dRFHG
BX#^1=O_G46c^a7A1:A,O6\<^e6_^N-d,0WU<5ENJ-L^9d9eH33/&]dQ&e]FGD87
Q-3c[5-2A<JFTdB9OVM,f>N0aNY#C5#+188&J5[N;e@gebY1GKZ,#f-(^+J@[&&#
.E-b&:/7b,7GHWgV\gH:S^O7Zd5@^1\FZ.Z65^2SOWJRB7&See;Gb9T>NTT40M5G
;;QJ8KJ)KK=@<#OK6-b_<a.GA&b3[.:;9I\3;_&K,L__A7@ZXP9@GcA:^F&.Q]IO
cO6;/D?P=+7JPD-RNY^6?f/P@PPNT8)L#O375YU6gN?W=Y#<_<_GZGgBR\N)B+ZO
VG25K<>/^2([+cS?+G)c1<.#EZAOVJ\CWgD[1O-1]SFAQSWK5aJ1=QN-.2]PL5PJ
+V(>P-cW:9N6MU1YC;,.4Vd_7E[WcTW/a(4XC/RBe]HM/NX_GJXDW/6eF-5@WF-,
ccTe[=2T@ZDLF&ZCE]fg&M;X?&gHO2XC>ANT=S,38OT;\?^bXV;5BcK-22W8>L^+
@JB=;AFOc^H^8@>E-E#aKJG]:eT+-W[T^F=KBNG\&KOSZ<dQfA\P+Y#Kd?gMPbcN
&EZ/cF2S1:JR37S:[Q=_;f@?<7WNbFf0@WL,6^gPK9[VbTGWUE;RC+J0BKY.2@)b
D+S6KKCN6#T3@+XM0g1:,U1JP-6&\eXY84_9;U5N:#ZcVFUcLTTMKN@3+dV(dD),
16W0K6;VDG<dgDZ??63:LbfJ_\J?1fc):9=ZKa-:C1=JJP2097E8T\;=EGKJM<HH
&UK6DZ@4QQ_8IX)ZY5A]APUJ:1F^2CBYa/YcKDM4N^HK8?)WS8\ETJ5+VB.G,]-a
MdfN446F1<1\b/<PJ8f0FBQE7F<)_NM9<H(P^69EbSS1AMYdSRa)6IU=/,9A<?_H
a?NAV^HIG.+d>d\4XYLEQWe@7YPfC>#L93J40V^^@&ARRD<^9>V_Rg.f-M9g8(Cd
[3T+#780-8)3VeZ#dNAD,Pf[.b92/fG+-.RfUB#V1(:\e;D[cNb^P8YLCVV-G57I
K^]^3K+/F3e-N8b/P6V70O5H]H4V7PC6_I)QEH#9Z,A(;Q/.c,L^fIc7D)WOdR0g
W6ST.#KY#eP>UA?aSMT2)C19D.>636EgNL-RN-8?b9IJe)P:3[1b#>a^CUYU.?:V
46QQ<CB3GC>63B-;O)NWFQf_Dc5E65W7(K.e#Z&<&cLA74:bX2<(O8d2M].[]^;7
63ef(/_M95_<&gH[;NJ_I&46N^#L[VJ_(?/b;._b[AG[a]]N;K@/6M5?\801HNgC
1CKOb69)9[&0/&=WSb8gfMdN1HgD^DW9R0J0K\5+9]OI+B-e^#4=cZYeS/d&081O
T33UA</R)e](VIL_5(K\+e>8^_e&:/]JIaGaO3BD]O;)8[\AR@YXP5cd&g#eDP,Y
,YP3#:Da&:W5KcXWD2a+cZESV-1C1HYf92EU<]0H9cZI,8/I.=0+A@R]+aFU#X5d
LXN-B4Q[R7^CJ.A/PXJ)MbG@UJT6EbB6OX8LX)B^7UPVcPc)<_U,A24C6KQU)<f1
gD,fF@^@b-+[dZDg.4)8BS;f4;]C];7ED3\RKc^AaaVT4Fg&<R0O.[V30V5QZ8B[
V<^R_Ka4KR\_QFH@LDLcM=KNdQ-UUE0Rd[CbUX(4Q#]9a.>@RV6C.755DeGUZ5;3
>[,f:aSa?\Q8/K<=.Q#HgED/+fbA;TA+OL9-XeP>E,9X23-R)@D&>RF-1G1d16Qe
KQ-<f>_M#)JH-c1(R8cL:+>@F\L^/\+T6V5<N<1S;.cQUL/F;E_4#4e:OVb[R13-
GMR[>4fM2>5dd8\3a_SgHcYS33g3ED;YN_Va,(e<>-L#A:b2d^[,YB+4X=Ag?==9
feVa&#DeH(152F:T9UMCS&GAH3<?5e4\I=UV]GOa:5M6,0g;/PXJ.1d5-A##DZKf
FGC&>N;X[23(?BP<RL;W;H1B\H3dN441C]Y]B=.eW1U)6I>8HK4=A-#KJG@1-+Ne
<TE:/NIJ0@RAX8)1c34W?,(g9[UM[GeadD^8E2[70=;/-WRKF-H20E]S#@UPNO-1
2Z6GO]g5:RGLNI6=YAO,^[<A=TNYNge@+4d6eP_+f_X7He)CQ?UX0,GTgO94T/,a
9NGI1BdPEe9NOC+;aG0?9X84;PWKD7\>3\c>3#10H)Y0@=HVO^]9Q6Z8HcT(H=KT
=G.4MOAc7K)U+G,O,eCTKFYF&S,;GF14WY1[(d>1a.30#DUK.,c2#Q3<aLSc;#M4
RN.3E07]-B>F#R@(cXE;F0KaBX9aOA)dP#8QO.T&:R=K[9K@1f-A/-AOBNg/&d#Y
f>@?8S>a]6U-9LAZaCX(2\X_FI>,8[,[b^:[ZKE@),gbG8<+8W9Gf&XK++15^)Z=
592O-84-_N/VGe5U46[G#Fa63JGRFKX3EF2.@EYY37A<#_T4@d@5HB/9/Jfb?a#X
DLJDD[)2&@b_RP7V5R6d.I)e(XP9&8^EBKN&fE;dP=ggeYc=T]@Fe/GPca/:6F#6
WM4=GY8+RE_:?g?/I1Ca:#A[_cJ=[AT:GW5]8bH(We9-9CHV?,dK/Z2BZS+NHK.P
\8;P.\4TBZ;:eLcCA_W1a5D-5_aORcXd8=be(_c\I@QEV6KMY0N]JJNV<6Vd3WH>
J2/X_@GaI4_W3FE2WVa-EH5_?^>5CE?30cCeV;DJ/.?9D[1[d<08;://C0UF3U80
5C3&6\:GK1#4AWOT9-aeP/CK[O;dN3,8fE614dTY\5;S=(DOg8)QbQD+Y3RU,5b6
9_#N5aVYB>&^,-?ffQY+gI6PP>5[6g4B[_/PN6I:]aMW5e3@W[T:0TH?_T>=6>_N
QSFJY,.)FN=6]:5:IdEXX=ES.CfZ;7\:#Y;3<[e#Ud5H##[cQ;T\L.T9ZA2\=<S)
.+Y+<O@@A7bR?ZT^T=2NJG(9^g&E;=1>0M[\6>JE<F5DHTVD1D.@8^#ICTe#2?Me
3AKA0^TG\._ReK0)DgW^OV0BFS_f,2AN@2G53K[UF&P6@>@XCJH=RBA1EP/9+dCU
YFaPbOD[1Z@K4QMZ7H2dZ#@3OS3A>3(+3OJc1^:=9YY35B@/RK=&K+R0c5e,CWFI
,B2d\<-VT4Z:<be<L:?5_N>;QC0>G\&=,_8CQ7[+/I;+/c.cGTNDY;gP4?@9Ma(9
gdK.g#Bf[e#018L/\Q1&,T+-E3PI36[#KV6>43B?4)8]dTL9,ZJ@?.I]];/K^##R
eB@SC]f<dIMLEeR-G5A0bZ0edOSB#@DDF4YZZY+BbI]N#3BXb=<.OBJ=dH?#UGPX
5VW.Z><FGYDMLX??HXc&B&ZVI3_XHRXE4Q:]OL=0>0K.,Z^\A&GL_,e^=@8^2L]g
,3SZ35K8GBUMF0UIJ(TY?YOR^IC?3=-XZ&@2KCCZ@T5\CN-0K]B7#;P;-[H??3(T
D<W^.E(?\7U^dK-3DOQEE6dP0T9^]ebQAL#W@L+355Z#7E^?OaWfM@QXD8<b2a5C
?,#A>L/UNG25,Y/T1-FJ)S]Q]^2[R>Z)?KG&XB.Sc:_:HcS8M]@Z&(CHJ0:PKEB4
;JfE#&/Y.Q1c1J#WA[YBf_ggR1<W&YPY;((<_bX?B<<QN<=,/TG1#8MKEAA<G.T7
8(E;RD,be:fT.7:7LH8M)SI7>_RY[[@AdAV&[dM[VV4BW1eL\@;7C^(OcS_C),])
1H+:2Me5c@/TO.7L7<^Db)N^ADW[P9V#DV6(+g.GbXb;H#H<c-IM@eU]8a.dFcA4
2Bc-B@BGb/EAg40c?^?A/,1A95=f-8^/=3YOD4TR2M2-aY=f#]Q>+Y+F(1(:K>+(
5XCH-I@BA0ggOVWQ_78g5Mc,W+TD\0b.GP/19U9,Q3E08]8=BVg,MHK@,-9RCYL]
^2M2&SgCXLA>B^aZQd5)X6+6K^#Y(/#+P82=W#3/Q.aIb40R;PJ,]&Ife=(=3KT-
aA_O=QLa3KeA3CAgT(Jb?]7S^e:R#K-Tde2[:,)]cLWVVHQC6Hb3Fa85UPgg(>Ff
a=^<99QR6)Z:M4I^_2@TH+&/=S/eI9A8O>P2V+<,(_,]Z;>EW1Q+b_RdMX9dS0A]
#e<-eF)A3abaP/<@X=../RZ2.B6KdAY[]E^JXf?gXK(.0WV,Q-g<N#_T]NG^)DYU
/Nc;XH4\V<c=R6B>8]<_cGZP;)R@,a.OaDf(;Q&;6c+eaN4AN<S7PU3bdL^J-1g#
QaQ7>S1@F-P.X377]SW#:.UVPbYa^f4DGZ:JFd+bcQg-OHcRgba?BTCKeD^F9BO.
(a/XPGF[eD3PE[-=3((OMeFb[?5H#(>EWGB^a8P7\RVEeb\-BPCT((0O1KP9+.=0
)AC<)<>\]BgZEEa_7U2IgPV(CgJ1B@+3;EOf-.Ue(YUHR#EQIa8H\5@MJ.ECbPU0
D^RGb2b:+CS>O(&,F9eF5M>[<I^c\Z(&G>Y@\LbBDd&SYH-+<J-;&&O]GRY01L0R
OEgOXUCR:+RJJH^QA?#0Bg709WdSI4O+?)f9f)ZRfG9abB>fTZdaD52G.C5UOe#Z
]\R7.PPV=AL+8^T,_[G8RT&R544/D]EPODEP6H_@+cM=Ia[F\V7\MY<?Rd??[\Se
[8O0<BMPf7=SaA\=FD?I.OgS.1U<I7Y,?U=8Wa?9,Y1:-YV_8\_=Cebf=\GO<2]^
F&><>5\[2,5Bd&fGb;RX1W8,=SOK(K2<<@eT/@#E2(2e(=0(Mf)SNM?M,LC?)\Kc
]3gWbSLK:?gO3/Q3\fG,/VJ=Y@ROe</B:cT#APS73[QEbZ_If5SIBOT53;C1>E(M
B&a:KZ-M4IHHRa]B6AMJ&6V:AB0X#8:?GA;-fNPR,0Y<Z+Oc0T)[MKS\[fQTf:bP
-[TB2T<GLNQ:_H91=?c7b^3)Z;V=DOdWABB/b<e,(@>#4.6)-?>c-(8S,8OXTc>1
ZB#Ta0FKOWNI7&<8aJ:QE54B^#3@U90C7QLJJ@PPT9#IA=c)dJ7Y12bDSWU\B)])
(1>I62J1#>8.d;Tb0ZJe?A<?T.EfRaDN#5LG[gDKT?)V:ed?WaHc6T/(^XT3\b5?
BY=W:,dRNQM4NX#QIU4P?#NJU=,AY#?0VbM=[@K#H])/#7HT5[O@>-=NQNU2<B=P
#&\YYCWV>,R70L(Tb0X.2R/EMLQ;0\#-MFX;7MJW?@&=3NMcMfZ5HV=/bRDEEWK&
30YU^[82\e\=38RRf[X?XEXVAa41@_5B+8)[0R>]\C]O0aENIA1HLXD?]8+P4V+;
R\?NC3Wf,QM[VH..fY];8=R:DZ@.?;\UL<FYHU>5HXf&eacNJ&=#e)Z9a^W1,_Id
N;EHb00I\RcAD2ZW:1DS^.^RK&@I3:]Tg8(O4>[SQOU_5YNJ7ELcPc[H]cSSLB.<
/#?1>DRgCNL/2^3.PTV+a9A#([FAgWOM/7W/1#H,YHRE0Q-Z/,<+=ZDbbOcH=##7
K+\NVL_<Pf54,Vc;c5Ob9JAbL=3b(-^(JAP8CM+c2b)f2D0297OAXgcRP(.(_]R/
e/N@U&I]O;8\T_KA1#CE/X)1#7@=EC2N26,_Z<ceUFe&bN+d4Y+COdE(-4<CK3X6
BVK>H7X7:;f\<;^9DO4Zb-SSc53(CUf^Dg5>gd>BRJgF7bJFY_g=<b^aPR8E)I[;
AAXb68Q0cP<3cRV7#N75GAg-#&(b/LT<J)Hb62ZV4N_E7aYC;@99D.X]J6MGgV:G
YL1K)[0.JZ@)XO<cSOfCfR63X\<A\-EP)5^SHM,b?Q&EX5:K4M;V37_WSQ0#?[Va
]MIS[J/ZHEZFZEZK1S&OD@fSb,-G=O:V;[[]6GB.+;^T<E#Y:/EBW#+A]V+@B+^3
G0WOY5QN4/Pb\X)1#ZB?<V5QfISI9O<H,#,=42,SH:A39VXPDWX41QMNX=(3a+Lf
PN8L^>_Z.HTU1EM87)gYEZ.(S4f)7S:B=[b:=-CIJZcB0UCAM80W3dQDL:E<D?-W
M5N3KfPY^<<>TURa6NA40883&R)Z@b/X2@-))(<#H2eZcW8eU<#&;#3d0.7)8D@<
AE_fTcd<6Q==OQEcY&S&29/L,;b12gEL,QHRN>Qe2ZLd:GJNK)7.SUP)#=bFIZK?
1G;_a:W4GHH5c:J;W=TH/K_+5Z=cJV@#HZ>-U]a2H=F,W,\_T3>CGUIJ4S\R7?aR
.H.&7g)ad<5E2)Yc^Bg9K@((Y9#A6]ZbG0_UXOI>-Zeb..:;.C@O/W)KbfL.HY<<
Q-VSXDYTZVR=a;N?:+&E]F3,JfQ+TT20=[&:OK_b3:f715R0YQ[A@6=c)G=1T@VO
GXcU)?S/.0_918d_RF=O@2]XT>?/5S._^\bW;X<BWaH9a6)DR,02HQ:.ET3/=cK4
B8aTNcN,WP5KGc[;9FJKO&ZY0-JeR0RYEO0^W0RESdOB:72P_VU4XQY))Z^[W_ab
82FADC;M8]MW\S).[<#Z:K\e6H>?O/#+0f)<QXfdM7bDB)dCH4]87ER5L),/)^SQ
SI?gNX86.Y3A-=0O.7BJcVKe2(c0<eXf#L3J-5#78KaFA5;MYY;ZG8GKd2)>G:W:
UgJCCPJH=L]2,<ZE1YHER7C[c>8WaaHC+9HEX.C?aMP/N[XK-(A#;L^7EF^T_AX:
eX?#55B9?AAfd:dM#QKeKBMW3=U1IBU_]/ZHI(TN1O/(d2X&fcd<K]DG8)R9R<(:
HW4-;A3_@&fH+L\?H?I\\^c_;?XX,1WBX0b/MV,MXGKC.W[9a4DdcUfISSP-JJAE
G9@4Q8[LMBAFS8EZ1^;aGQV&,#9(_JHX+S/gSRCC@[LIYP)>SN3fP\#;#gFE)-&3
3R34S=bQSB(66Q?NUNEB3eQTC:/&DK>/;57a:MVQIc=M:gg6O[2EF[X?Oca6C7b5
ZS?5\A4R)Z@0Cf7c@G\[\Q-R[&-1YH+OA:98:U)=9N=g7BdR_1.Y&2CM/[.e3c.#
#D-XdXCZ=4SQ(NfSJQ^O&6(Z?1:0HR5JbYb:<0EGAE>>5M\(,NA\-]YNF7a]VcLF
f3eQ<7<3c?N7(,F28GL19N;dO=\X[9#/&KV&?TR8)OXJI/bN/[5>@M@&a.7Y2__X
9T.;aWB@QFEa2P(^g+Y,=NLXA5e#BP>Q_Oa_d^/^HJG]&?EC>THA9=/c#cI,(dNK
O^;aQg9;(?D.(N22R<YSC(Ee:MIZecgdT)cML(G_WTRV\BJ2>YAZYCTC];GYO<+b
=+U?e#[E,45:GNcHO:1:P)RR>1GN)FR=]1ZM^g91-Z1265&)]L32Z5:#gD8)L.gI
U96_1[Q<c#LQa.8<PZJ/4#W#G#JU\:ZYgX>FP:<Y]DabeYA:gG+5^F>KZE;C8FX^
gICHd.H<4A[CAKe_KZ.g\GT(N@=LW[53S0S(XXIWXG7f4<AX8aaU=S/9J/J)&OXG
(_c&FQ^F,Y+abPeOSC?2:^R_JadGMb]fE7g]V@(=dc(+:-c8.(/I]AF&5-M8U6F.
5?aA)]K39AJ9,deU(G>&\#/DZBe#aGYDUH2:;,ScR+639:a5-4+__D8DIDJW?-P=
Z[2?_^<IFM6R/[K,-?N;c4GVAXJSD:Mda_J6H81FgA\eVVc/E,MSA+2-H9MDd\[2
YDY+(c^_+D@b7<=R(:4//;eQH)0.d?@+cf.RVAFZ?^?,fH52^J3\GaaWRL+)H\FX
W)3[G/44aTf(g5+cLXEL1=>dD:=bQ+d>?[-P,L#C,.]+\-BKQ+(>+,-dgUJW[+@5
.LH^b#WT+dZ\+2R1,H9XOQY_BQOg3&A+bTeP_V0]IH/+5Pf:KX&cJ<RPL?X#(eR@
YQ>H-FgD9D+;UD[<_/aQVWa12E6EfTbHYc]g3+80_X[9Qg=<@;_Q;cWaS-(aHPW]
),Z,)YbPJeHUXe7@\9Pg)g;6/E5KAe2&aUBc43K3/=M4^RS-f:;O_L,8F>#gdX^K
9^]Cc8FJeNIA&OC2JgYL@O9H78(DN7UM/8[V_+2If_;2dfXF]HafLY(DgQ=gPHAF
S^17L2+=JE&IARR@?c:NT)UfTGafD1\ZJ7@b,B(X()W]>_2eZKPfLW=YGPPT]Vag
,#E00ATU1D^KVa0N]&RFV2[,H0V.bN,ceL\bTKCPeJ(X_OE_++\=6[@3QIgNb,Fc
HW9>0_a6S:/dQS)0DDW[B8#e[B8]0CJ>/J0.:9DVLVEG(U:_ef+R4N@W8c,81<V>
028GW<[#c@_C:_OD-g2YgZe,@X)OgB>+J->0.>?H2MVVH>gg<<Sa(P6X-L</F3LC
P\92-@^=@]2f#@F;#SC38]L0MTDE:PUZMSMZ@?-L8S-RcTD<N&3?K8\@:NaH?aF3
XOYJO<\@+;IW-Ye&aV,Yf23PVa.>3SWWe?#SgZAN?_BW6e9X&Ygf+X>O,Z)6^8AJ
0E:C+8W\0(a1PcWM7MR<gRP+=bRX=@]U=b7:3K,&=K?=EV]-C3+_WD2]6UG<)e\:
TAcCPQ9E]7YZ,-DC.Z+,M>[&A4)@2GY@Y/HeR>X85L>b\QYV>0Af.Q^aF7/,>V:5
NgBDD85L&.R<LM78]UCE8NScf9I+5RX^C&=<g3G\Ce7;4>Pb9f+M\\-g/QQ9J+?M
aQH-RCZD=PU@A_RH2)<QV),5]RGb9B@ID66@XG6QV_V/1g25;O@3P7_SGA3E@EVR
W^J@A5XfGN)gP-@c+8RLMM(+U)-KN\Q.GEX^P.e8]g=?9WI7&9ecTNR]XF5Z?;)=
OZ8ZP_M[-W)aQ)>0S9)=W0Y.C&GEBO-cB3c&;V.KLccR/4KN]]IX20cW[T)#DdMD
D[UL8O6VOf:Q\T(_)f?c5JUQIB4YAT?G</.F4>1NKHbbc-4E<==_0H;BQ(175QPZ
[5<67M.a\9[9+_9-O1b2V737HH#96Fd<1Q0Y62/0>U-Ea8SB_=9,YQEMW+4a3P:F
LT-FQU:.g2Vb3E?\0&1LZ99^B8N-Wb(IDH&[\@LE:U[IIB4;L>/M=F@Z;7ZId/,c
#V7((ZA3e4Z>1T?W0Mg^ee#Xa.=):[\MbJE+@=Y?QYI?86Q+58OJ(=K(L[FS7W1U
6ET^)d0SfC^\7f/[A=XX->SP>>:9QO#SfW==:K_7<0)906R871Jc5R7)e-O-;Va9
S>8a99T>Ja79a#)Z\.:B#]F7Be)EeJ1(]_YR5Y>ONP52KEa3c@:;1U1DOSP9fT8,
Qbg//_#\,7ccc(:OaRG6\XXe7gQWUO9]IG(U,XR7:5BAd+@]P/O4J53495KaRKG6
UTY,bO(GbG2L/+-QFg(E)bO,W#D-[CX?=:/2[+:)^9SLF)X),+d=-W7O<G&LM9;9
Z+-Y(bV:L6->G@2.\XOMb]1+_=&(,+W=IM^ed81)QSbA0-J=H+3>?S>2TAJ#7WT\
:1Af&ALMY1O=<580,@(7WB:@f_eT#B)NSb?cWWB2^(S.&dMXAFW;-A-T;/:X@.XQ
<ce8?V6.DPE)Od\>#U62LNP56B6Rc_2))FcRJ353K#.IE>:;?^-.]DfYAO]ZIF,B
HGKYT5\B4GC--TG:AA]5C(c.M\_FV9=gAT6Y#3D\He8HOS@?(EJ=X.YSX+EMQ?eC
>9_+c-C+H4)=IeGM648]@SU_8BE/Z]&+B1LM9g6NT#9cW1eE8.CPAS?M3H^2GR\X
_EMXf2c+G7R&@8K9B3Lg?9aH+H0MdDRRFe#X5TCH,(f&6&_,\T7?Y4-#_WD\>I<d
cRU_P>?@58,1Z/K-D3aQ=:Rb@d3Z)M-QVF8-DC_4ff:(/NMX#;A.AUL;d498&:C1
.\75T.T30SJ8OH@ZXI#S8\1&9M;WH7YbQSA&70Ac;]503dZO@4I/N#d3_IdR1K_c
52bbV]^#0Y;@f:#;J=B1/MW)0,g_IYJ)6b^GEW6B#9W\U6bb2HgJC_KBcE;E]T#1
d8cf/7-+WV6=F^-da\I?XH;(Z]bHgIOZc^dDTK&,?KCdNE=8ELM<4/45Ve=J7[@3
0OI4A&NBfYA2HGH6De&.5g0GTS>R-c=4<c^AM2a;f-QK]3U_O-)Z&X7PV-T\0Ka#
.++d+#I]YYH=+1R4+=GHY6)FDg\9TTF3_FS-V6/USN8OeZBVGRf>Vg9H3V(A@)cG
^WO&L6[4.cTb@/JWY=-DD1-e0<0)E88IPAec/O)=T7#HG=Z^GL<0Gac4;4XBFRc:
HTMFA&#eTYEF-<&Wg[bXOIaZYY[5RWL)<b.8HQ&gQPUM0a6MX4+OID/?ZPU\+C/?
e3W-P1N^.8+OP2f)=]EeL4V_F_]?/H?)&QU\HQIfKIT@K@T,GH2O9_3+YS9>1M86
(OX0AKE@(g8RR/_bGe\<+U^FdaULMbV/aE[9/+\f@S56a=?O\&FOW=^b]B2D+>Dg
K=cZL/a.Q75H?]cF[8/I\DYWT1J&_CIgP=P_#EdO+B:MKeGW=TD=Z2Zc.;XR,8B9
=]gecE7)-F+<J=VG36KP0:B26OdBH3aKG9TM(EC@&G=<>:Z/6_3T)0:KYI5/:R,M
8Z=f,@)UW)24WbK0:X:N]XHbe;IQHW7MA^Jg]bX0G=\b4af43OZ#KPVE742T0EW-
.@OJP.;=(T(BY\:#R]3;W[6QR0+U=>3^GP2Y#4(3\c)3g&.Ide1+/[UDE;[f;f.#
BPPC>8IJN9Y;9VMUUY:6\eO,J+2LM+-JX3/,J#&@J=\,089OZ9.XWY/20KB)YDD\
.C6P,3B1\S6@K@\-LFD7_,;-E:7@RI[AXZ@&1\R3:;P>H,=KLJW4JZ4Ug=?_USDT
4T)@A9ROP7^D&MWX89W\9)0HIXX6f,4N_b;BD6E@LA;R==aXZ>1Q=.5I?Qed-?<-
#=Z&]9X:]BPg7E@U;XJR98+e\?;P8Y\ZeA\]J70KR6\(-#7VX=IJ:0K&VI&=eV]]
HI(H&;beQ14eT7S6WW/97?+N;bEcG4Q11g_0SEP@S+Q5g:@Jd]-f1/X>WH80gH]O
CD\J73=O]W[U\;_]5LWfe1\SKc#,6#3K+>[/=ED@2f<A)#UKQ(DVgCLGOUR8MSJR
((?<N3\\8C5d)S+3+.T.W=NRLKAYP<G\0C:^#0b&[W&6+:ESS^2TK6RM)OeJ0]AC
UR55,4Z+EegRZOFS?Z-.S[Z:;)DEP\ff:K+-b7AYW])N5#3dWVLNB^e)TQ0;HOdB
\[O/-F\5-7DKJ+3M4d+@@KG\Sbb,0-?@ES&dZ9)>K7\_(;MeQ_TC+OTH:VDN,6E)
[BfRdLV];C\XFffJI/<IB5>_B2NE>7U-KC\Og)<?Ff3XMG;Wb++0<a\=eg:YF[ZZ
^NFUS7JfFgaIfK8Fg[_L6aX=X?ILJ:eM)NO.VeGe>?d\Y[MFV=8)R18YJ>5c9BU4
?]dJ;^.c]bR+B]9/L=gYV9]>6Ma0PcL;?1^Ecb+.f-CJbG7B&C(:1?-a&d]9HDOJ
fdNVR-Z8WIBS)]_,H?7#:=W_6XJ];)<Q9NQ/2F-LL<&LTG],HdUN3;RFgJ#Ab-#?
FZb[2;DTVNQ?5@X1+M@#;HDHZ7dTf<QL+^B\:@?5Ng\=Q.PK8)D,?eOeQ1eR+cZT
EG#+-[aX[^;@f.PA&^Q8\V^)<#Z<Ag-b6^@5J3D<WC@)B=O@NQPRE.:N(.R?KK&8
8a&+L1d]JV]K,06MS=NaGT-:[c2f;W6:?T=W#W/0=MSBaCYUC@?UG3I\7bg4N^Z^
L(ZCf4#S5g-R7S&92@VWd_dIAHY\Pd]de7,MTH:MD+DU]Fb#88IBCe:#g2.=O+a?
U\TTN)5WdGD_e<I@)Jd?0C_ISGd:MF[#HP@>RW<DTAe&Be4ZeNZC.0BU&YCSce-2
F#-C+XHZIcO>/U>D[:GB5G9OP8dg3d^[7^)]SA:;CMBF5^DC2>L?:fAa5-8-f;D+
-/AF]RGNWG9[F@YNX\G=-_23MN7,TH,4U([-]=;BS/=]&7L(J1AeX0Fb\a-<.UTY
1>KN&):@6c)+4Y9#,.0B>.)+06_CegY,WCec?/\3.aNbO1dcAV;(b2C5eRLN&B<V
UG9<8:TPL7@AZ/4e(P852U@]9+39SfTD_JJG]RLHSNZOJ3@cEJ]A+?GW=[)YA/JT
BHR?d\VS\69;&Q1#QX^HCK]0a&7(<gFJbZYCQ+6ZK,H=40CER^@7a3GP//()A@AS
\c[H;N)VJBQ_?cYfOQ>H/+&1fb.R-EPXBDBW,=A4(^M&M(AI3BL8+I,Zd^1VP&a>
5+G)JU1VfH;1=^NDJFR-1G?23XQ-[-)P#SKRBfe=]5[;9IB=Gg@97a=F#&:D9YaP
(_#@KHHSAbZ4<D?P=f22-&M:-.Nf:T):&VY-TO?2P,RgYI^9B7<=?Af3\->W7UM(
>]1bG)P[Z]JM-aWKfY/c++E.>I<(d:cP)AR+@R97Tfd&?1AaJ=8&=(2(A:G92[Nf
1&N/M[b30M@e\W[MWg4Q_\GGgW4S?0-eSb:&VBNM2F6&#LO.#;17\39-GJP.>1._
d50XO5Ia:CWP>55[g(bAcZ_\[?P9O8F=&B[b1&bK=dG3F>+G5b\+cE>EA@S?]-WS
)#8A#)=];)Rcd0S@^.#c)a[b<H-])3PVH=>K1OB(RcaafQ31CA&VD3,DcIR8E:[c
Hb[M(J6/43QCQ#@3ggZ;Q&([;][YAWZCH5N/;>62#[e)D5+DQ&OVC_]g(\]PNDF9
EFABGMbYV<WFJT;I?G0O2&VWaY#8XcHf@E5<UKdXJfe\_gFSPSR2P/>4;9Z+:S+J
O28VC+I1OBD9F\Y1.UE>D@4a;BJTP6.NI^,Q-_d.HIcAfL^=\]@fOFf>&=7#_:S>
c[WOf,5Of:S_9]V..)#B&V_8)/Y0,5V;F^T@R2Ia^I/]_:Z<X&[b14U64;8>=\]6
6SKN+Sf7908g_FII+E/\b8:5IbM/K=^6_a?V19^]>R^&cKQ-BVZOIH^4S(6/JQSX
<T<VVBQHUE5BX@E^:^VH4/>3<Vc47,ZEA0XK]&ZXG(@4#a9WSWWUDW&9-df)>20g
)]8#Z[fX)#SR:]>\XK.VcZGF]c-OM=QKQ@P1W/4.YL5J@?U]68Y#XOQ18<2VN+2X
_+7BadUBD-X:L#G&6Q,@3RHe-DCZ33KADU1XX07;B_f^6/)HbJ[JLX=C6<\_-1O+
G4I]/E)\PL-H&>XTEJ5ZD1#2.<3W=W9:d--P)HU8:GN.fIZ-<#gaCES<GD1[+(G)
Bc&8H4IdGDWM\c?Y;7T?HA1>I<?1K;,VL)HDNWJGDf[7M?2-B:E2/eS2_-A/&Fc>
;aK]Ha)XU=3IT#3?OPQV0R/F[S3+Z=K@.Va17>:]WQM3?(/<G,OQ0FBA_cUU<?Wa
;THHGAHECcIO/9a#aV)UK2J@;:M57?UDOJ(0Dcb7LeH-/[P[9;>YH+\3P:HK)g=K
Qb.:);IMDg319PgdN.SOf.9IMN(CS;R6[Bc=cg\-OV:Z9UHS.Bg:ZeO0-85/484U
ZUC/(^L?g@GF67D0MOT@aL&_I0gEBg&>;Q@,(JbdF]E?N(\E#SQS?1X_&#?R]>)U
&<AJ7JS^BWJe5Oe@92SJ/CS<OPf>#^&P&<,MQB]N[D#S7LA]N1Y.\ZPW4J)9cH)g
^A9;RM]SI2L&94::eXURd+B\b0>])2729M<a/V4_cXG3,e6POFVD7>H-GG&2.5T_
eU]QE,]ZXfYNZ(DM#0KD48FE=>XNf<UdJD^_2Q1QWbM#__LM;QW3IfE0Ia/AUZM_
<21UFc^-6:XT:Vg7gJ4X[KC2GU0@[6XU)PY/.1^a]HJXPKFaF?I+@>=DMOWBS;YJ
e)V0TSC9PP/X-L-(UdU95A?<\[BJJ^4WQJ@;?f;BeET<B;#f2D.Q+g0Be2_D([c;
C/OFGb.LJT&I[>,]5a^(]9+=32\<1)YRc5@<WS8O\H-4/>^<C\\7WMCRMP=238WX
<fC_RV3D76>b[?Z#=b+)b?>Ue7SXI9#O6M\H&Q^KX#G58DVVT;1&[CeBO70g8Z@Q
Ocb:S;28_EN+gHXK[4FHGM?C+^.^<56:9<4@OT[&a^DfeWaZ],6>T\/0BEMHT?R_
RLc8HK3=ZPU#ZdOFZ:\S3^+c,67(AfD(f^aW-gA7_U)PJcJE,2JD92e<Q_^3fN_1
1(5d?.DTX^Y,]Q#WWIY<F5E419GA?1>DZYN0,OTbF1SRN(][35XVNP\(cS\,_V03
L;\G7A(BAE:]-;2;T+.1.O[.TFL3JQDO(I7XZ0<T[LfOL,0fN\FIQYG#+3b\S=+?
.a,fLFY:0C(d=BK^P>3PAG?_eL]eG3N.@;S<8Q:PGD-68_:CZR6AM=\[+fK&<e6N
PL@95RfKeI7#1f\H.9@2\.WEILa5<^bQ-7KME,/=9gbCHXMcHAB5A.e5TA<be\5K
If=KcF#.-&)E<)XLeFBd\2EF3,6@)\=UYPGLFD9QP<\#\G8984DEH1#+3U\5>WgT
CJCV#V&aVBg#<.2I^3)87B+2EU/</_+XNFPd\9Y@I#77[J>KgH<ecJU?Hg+BY8&T
-@PPRU+ce^R/aHXL.>+TFL.[,.]HD?CF[IPITf^\eg3_HgH=A&#);EbP9WC)D>c+
bU8X(]A40<]GM0BG;#[8HFY8^&IT]Xd#RC&6aS88;54fN^9@<76XB:Y;M=6X/&C>
>4cf83aQgTH:YP0FM^=a_FJ3+Y^T8gIT;d#9/V27Ba\&f+3G/9&&OcK#28[;g(08
(0AJZPGdSHC@Mg(Oe[abSfbPb)HC2PdZ9dIY2E>:R7>>)2+#e5FP;Qb<Z[HJMfV)
3JESOP45<-Q9=aR?X/G&77,d.QRe?/>/gB,AbG1F9Y.2a;]PFHY:S7bT>6.2HQMb
g=RWJ19RaR,KGae@]&PL/DWQD8N16PfXK.IA^g_g_??b7ZIC-.bD>3X/QaV=?d(Y
BPH8T-RNV017T76Pc.U9eG^2)(?.EcSd>eF>=1TEBaf_41^C>88),BJ;P(5H(#LQ
,3-?T7F7f;.QZcdD)5.<R-?/8/U-Hg?G&.\M8:a+(NCY.7I)G0LNFG/(N@@]Z9SF
87-:\:.1U(L[4,^>8<Yc7>OJLP:<#e@KG4SG0)Na/P7/7b3S+40Ca(VB6AGaO1JR
b\C\0Db]H>:a-T=fdBE?P@2E@O.=/VHG7?3?,DLV7;FR=P6KJ@FJM,MSH?WFEXM0
&/7K<XV\A&[G6]-Q(dXd36S1e>Q<>/M/Z=8R/e-SX#SD@2V.,fFX^/@C=,bXQ=RE
Y()G_8KP<Kb#>T_RH6\Y?JWbO0Uag3S3._Q1HS/2E&(S&89&RLZ)Vc6ADTY1.XYK
@SV56?ag]9B/3H=bGJ)YSgYKHVO-ffS9U+@=4Rf:QcW_B^?E=R=W=@?O#@GL.B1-
0:7XKQV+XaWI9P<XeZ(0gIH.(:YPNX0c^B\ePZ7S,>9UgGKa4=DfXW2KE@,82<f[
D;ccJD1#@GT>S:73YJ++G<3D3bYFG#A5I2Wg3E-<R)A?>5/Oe&9XV?:cCg(&,_:K
UC5@W&7FEb-JLW@:59&>8]f4-N54;FTHPdYOSOc7gF_(1f+G<HbPB0-+e7/N#Za8
c0I6LW>MG2.M]_LcIHL@E3>ZY9Y,gAX;#2^WNaA(]P=L3)4[KBbNC[b&V[1@d[?F
W_R-=2P@<6P=Sg_3#M=;:IAO+=PQ\2W.cB&8U)+3eKB6QP0eeC>+LXFQ5511<Q3^
=O=_DKf&F3c^>+_:FED[-B-8@6-.XR-J#V^6F;f6G_;48OB&V24YT+cUMN@ZKMJB
Y.:3?IX,#YWK><4QDEe7[HJ2BK-7Q:MRecVE#7JSWWFBC6=@W4O-LOc\))BXLP>O
+3N#K8<P-YRX<I,17B<<\L+?VC0DM5SaDTBWEf\&LOS3W=gHRM/:bfR<cbd2-3WB
MFM->8;FVTUJ)Vf,7Z[CX>&;3BZ_e=IZHZ(?B1-;DSb7Y\&L7Y4];??O6+GWQ;O-
+F31[<1TJ-:Da?&0KVU:Y>B]38&a/EA[XL2Ge\I>G^Z#=F)DEJ>V.P#L,\9)N^W8
]#L(B8SZ?HNE[T,_N,NDb4Eb[KAGe?14HS908D\/NFH91:Vb?-T_E0+I_XFS(fYL
L:89(6CXKUL,>.C(CRVW;>)3[6B(7&0BG77TP75RMD>_4e03FWT(Ef\EOdZ>ETBM
A#IVJV5K-d=ISa=X<07,ec8(J7gI_<2(cEDHN0?FS/NDS:GNC7J4WSN1#a\==e6:
AGV<Y>GbHB&fJ&_7=#S#;6@0^M5\;eg4EP8SP_-.eHcVDU#Zf^_(K,DeASEc.PY)
:SV]Y)_[OJa.^)eATUC_e3bMbg]_Qc0<&094KT@WTV?2863Pd]1aEaDBDE,WCAJ2
_[>128DXI,C(e2dd#JHUPPZ>]LK4:Lb<(\#BD5X/?\>\DAX1?PH1.W<0K:XT7cY6
7YYS94=4ODXVQ3da/<-MX6AdSF^U^#g79F&Q+[VFg0MP(0c2V3/4fcF)5Qb^3+d@
@5eN,-D.+]aP.S28&,A8H(>DIg:G]DBB..&\+UOcE6DM5<C&J:JW,0@&YFJZ3Og[
MAcM0IFC8gGQR),R-P<;Md3@KFdS:@1DN:0YP_aJ39WURA[c>1JP/MJ<9:?7M5NK
DK3DZQ)g?2^R)R3_9=&<0566W+-gYV7d8ZMVc&c.DPVS-23g^9RK4;RD&>H7N.H,
MO>0SER=8WHXDe,TEW8GCG@8/8+BOAZ_XKM2D@8=eYeH#AbdT#9PKP_RZ5ZG9Q,H
P\(0W4:FD.2SO=^CHQ^BZY6-VA=d[P25SG1(NBCEJ3F=\02@9/JJ)eOddBRTSNLE
D0_YO\\FRBVPQI@\<W>\;\Tb?gJ[46c1(&EDGI<UZ=L.<K=Fa2g,YUVA57Yc,EaG
3^,6TB(8X+&FZY1CgEI,_Z__d?_X9R]P:Xg-aG=#K&9/f1fQ:-W>E307H/6<7@/a
9WE.+DCbTWDIcd7?<;0<Tb<6TU_PZIHMLUV^[gRg0LD^\(^a2Rf-UC5TG6>O+29e
RAKc6Wg,#V#@VdHV1UYY:61g+3BO^<?NRG9)RMXEJ5N;A1PSgL/NdCb<^:RIVI4K
aF(cfQc2WG1[NZ9#Rab0T_/caDERMS6dI[-P@^XR[VP1JS1UU?A_/QAEM)),,B_M
+)_a+DGK-<JITLXM=P#D3DMa2)KF^?&4WU2d@)5Z+(M.=XPD:.gcf,?Q+B:\b=gT
Z?EdGfS9&6(Z1@KJ=0#XaK[??f352K\OVMTKZ=dT[<NL>YO4Sdc<J5WZX=-7)FT/
C+1@a^dT^^f\_Zd[C0,WPL2[F))(Cb;?4aBWU\X5+_#SFX9SE1Kd[eH5>Nf219-P
EHg-c1<GG895>;0S+#SbgeaOMLP36DHcD-(;f>SP+4M8#;;5UXHG=>aBJ(VU3263
>EUQC:2&Q#f+#3cGZU7Bb0,Wc4+KdY7?^V(:[P@QPEEB/->D[)@9M?4b\5JYN9SR
PE[-^cee+WgGN/OL;X\?1V4_V=/+\eXD&[4/Y-1YAg-)9T6H)?]A_.<T@-3?<+8U
3eaC8A8/bPQQgN3R)B1E9(Z5@c3LXXR1cP7R^&BQE2UL+>KAS8K?XC8=5M:11eHb
^/>.K[CgFM?aO=17&&,X/&1Z6XP,b[_+Ye)J+,(8DZO55@0:3/8dA4<V2LJ<J8D=
cY=7WUH>Q;649aaWVWQe=(Je-,^=(Y[[M+9,4_V]A@[.TdV.YaW4#9SXZX<d[H<e
a5A?b<<;BW0N4R1TA3/fOCA&+1W9G#D.G.-?W]NcE@1PF5.I4VM4eZ9=MS:;R>5F
\SBC=(FD>V<gXYfT#VP#QN1N-(#,4?4818U<=W<6aBQ&JA79?FBRgGUIcAYXZa-Z
/M.af3G\FT1.?-R^=RS#?^a09V@466&&@W-b&LOHU;dfb>T>Y65(f4CTACQ;Ha&,
G);0#+,SHPGSD6^O0(9BOQ,8K=]J?S8()]VAcK=P;2f35J6FU^b9YN6-LZ\QT4X+
4Mf=NJ6Yf\JNE#G>(4>,52G[A4gXa.]UR9I^84gXcEUN]@)O;N]H5>7\/;bJa@d^
U2)BW:\6(<8f1GXNX#6SY/:Fa02QH?ZXN>6D@NUI-Qg_V(G/>Mb:0:I4[=U]?2&[
1R2.><9R\M/Jb9V90G=E\,2NR,Xc?46/gC;bU6#V--<#Kc^0V#7?D4439LX[AM+5
&S,EVXTCF&VU/>Lf/(R5E;:[Gc&M?0C6gIJaDAHZc^b\/19/AE[&C:5P(S2PX6DV
6D._XLYID&f?.E#<OZW,9P&UQSAIKcI>/cB?C_/;d[L6<.K@G?2GXZ)LUaTKa?IL
H.P&cDb;0c=GS\^gSJd48QGMP#U<Z7=FX@aK1IbLf@H&T+(UCHKMBNNXL8R@>^G,
LJLLROR1F,A1#SPF/2f-+UH\,UOUFSD5.f^R/->d+5=FS>Y[<c.g/X-YA@Q,QM@Q
2?ZIH@-V<=+e_g.G7fd5T\C)22(WS?bM<de8(bS8Pe_d1G/eWa8/IF;Red<UX#ZZ
Z)Y-NF(0Z(S#FB+d5f7H-F-81^2;>-0\RD1FE=59DYW9bT,5:KW2M]<ff_,B7a?e
AGXPcfae#5a216f#BBTUIQEUWa.]?>8a)W7&C5>1_YU:WV.@Z+5^Qg+E_agX8@:V
[P)I>F>eBY@\[Z<<_=YWIIW&M[;-.LIN5\Z2XQ=9b7CTI/#5-LW>Q?K;(+,J1+1&
F>,IQf/g>dVL/S7D&eM7+>V9^f,S7N;OMOH7D@c/+4D<R^E\Ec@F1)O)F)TT-X0S
9684NMbXC=SBGPU)fAL25=>bHR+3af=R0?O(@0^GJf1U^-SKY:egb_>ZAD.?8E@S
8NLA8JDLDN^Y6IeRN=XTgO=^]JgO(L?+I>C^-HgY^))7_\W_83@^>95\U,\VRRKb
#V_Qc.&L<,-5b:FU]BPff>Kg7d;P[>66G&EQTYW)6.EEPQLM]=+7BCc1\1)#K3Z^
&874IW8Q[a?W7&I@5GX^SF_4::7TGF@3A^EN:,RRKF>)PX&MV>WA@WPNQH<)Eg4L
.HHANXM+SeG)dJ6C(>?:F+B[HEB0eGd5LKU<7Z)\bS93dI8E^I1KD:M3?)?Z_F8W
J^9B16bP:_=K>f,ae>[_fT//MM=CG5W(VPS/M1#=XJK-U51R#I]/gaPf0RT&8MB6
4H?=HO39^g07YI/g-caT^-Hd>fF7N4B/819==V8M/L1D]CXc2<B6Ed/,>(.60cIg
[P469NG)3HKS)[?]Fg\</6&:30d7H/M+M<6,=4?UAP)UB-]XP5(=UQ+fKC&+L8X7
4@PP07([&+L#d_aU8CEL3dZ]><L6,1O&G)Y+PA]&OBe3^O(IHKDXg:/[ICPV>E-4
.cU4VVQ4(:?YcRHa@43+[a6P6BC0M[e5Kg5NHg2)Z[F>_bWg^c<Od^\Gd=YfO&9X
[-?\DBa2Hf(Ud(U^9,XU?ETB4+N,@IC-f]3e1CTE3P[V7Y.IT9MD)O>2dO0D4;7d
bD^DGW?8;HN2:DYE],7?BVEJ+KFVgd49;6EEC[N=/JK\/cHCCE&\A3[CG3O9B[[J
&L_[:\,IS8,&fK7Lad\c(AG\63IcMY8&@P>/@T,XXZXc?,JI[S=T525A8WHHFN[Y
cabd\P^c62S39TC;;Od6Cc>QS?3]5L#T+/C8^c^@KM)#<PMbfeQP67/J\9V<4VRL
GNS>)&O1//4[+e5TU=PX?G89bWGKV(e:YdDAS)_fUFG[.]Dg67.OGd#Q9D^Zf_LT
PJT/;P(\WIKPF6Aa^FU\[O[<]0.,.PLR0\L;c>A#Y_:b0-AVXBg2#3])_93Q4M.?
[:.+(b<bYEe:QC.YA/J_PM+Ba,YbEK/>&XLb36@dS@M98N::+1Xdff<5GGW#YSVM
@-Z(0S5c-7>).#KD:NRENI6>ad/_1EM94X+Ig?MV<-e_53D74a@]bYMDgQX?cPV;
_)V[YV<AL65_5IAGAe,4/MfHOd23]PVD6?X[>,eQUGd/FKcRdC.Ub3HIZR@]6a6V
^Z/-_YF<VG_-[25A\B-(;-MJC2C]:eLOMRQOL8WJWH3WbRU6FE=,LeU0A]OT)S#A
ZA8Ba&5.03_L(22f<3/?.X(L.GTdM09Y;0d()QbFYC5?]f]X:(;]I:G-S>[0DbE(
^U^Q7Rf6=<)0-<J<:=0aS\?\YH(N<RT)KR2BQJS3KeE=^Q\7B&aWI]..^.N.gHV>
-N;]HD#E@WH#4Ob1Y25UETU#:cL/Y>1_D60G7N/FNcIcVUMZ/L<J&-//E9.c90C<
?^J/?U>EPNCQbM;ZQb-c+5TA=W.&<<(J>d1gG81XB6;J27@CXU#EF>+LW](Ee2YL
X&8-NS^53Y&NO)=##@TG)8AcXI44?c[;&D^9MMMSCE3;?YR@D&:6J,Y.SL^&750e
XbI7\:TXT-dc;2</)[LQPcT#QC?,<],AZ6DSd4.+fUb+bSK,,^0;I:>I4XgI=N7\
XfCCW^a9d,@Q)3L&ROXZ=ILW=5c8P>NE9M@_GX^XgNBAc\PfYL7[9LW[^F2I:3F9
JF^b\BO6,ZG?V/aRVZb@;\1FNa3H@:cY6Rd:O);Ia#X69[569Bg5ED@+>]QZLHTd
?KRU(PaB/^Q30@?2&8A9fBWEeANGAF;&TEC\QH7YGDAXSf.5X+>6WOcbW#C3LdJP
[?.[[[gL#4242/eC\gfI,-8/8KR+MLKE#0:&+JOL:EW(NZ4,Z7SEWGDMFR+C7(@O
(4fM5K_(1d>I\TS:4OJM8OIL/W9H9XKT#>c)gH8CV^Q?f_f<I+2TH/;,]4We577e
1^VMJYXfJVO7H,@VaPZ_)6e/E(8L(D_BgO6PXQC002DWaC9LV2aN)@P6XF>IHdLf
4OS3);=b)gFO5[^@8VI8JQ9f?g4N47V15YDF2;BJQO=LE&ff?I/OgY]2Id4^UNX&
Uc+[HOVI@@K)T(BP<TW-VGT7TSNC+eASH?-98Q@5V+Za#0)?-f__a=3,D0eT2F=]
\TbWX@EK_,fAWC>OG/GLWeB#,]C5?G,9P8;IKFfPE(/\R=fJYCYOLA4cBcB/IP^.
NB].G3:=ZFcN8g&H?R.;_LK:F(/dPU[H?A[>RZ>>JBWDM4\cGL;f0.BFd>P<HY/Q
fLL;8;(Vd8Ob8USOO+()OfWL&4;2QL+B:FgO<=aP\b\#;dg<>DT-_;aZbe,92OVU
#H9)0c6T2/<dIDcF_Ad_]f\Y;6;PfDVKNHGQ8&+@/E@bFT\E;a=.B0W)/g3b]a\^
?G6496a/BI^?O4C_?JSQ2gH\WSDdX6A^WCG),62bC=dLEae6;?J/K.7-B1#5A?T3
#>UT1KMd<?LAGW4Hf27/R,c18abP55[FF5OZdfUB8DD>g([8\@8=5Og&-;H(?F_e
IN3dL&dFKL_NH(2L#a;LOEFHXEeeM4<gRG8<3CJ8+^99,6\0H\XZXFNcDJ=WRRTT
KdEQ;e-RI\:g](ODYSB8Y5&<+:_4,b>H]5->[>[Y2aLA-9a?ZEC=8[XFaQbP&P9&
?4CUIW/X:PeT9[@g[]9:C=\((D:]_->RQ[H^9;-gU2?27-Z-;T62.1US&2;e#^II
f.#M8Y[a,]RG0/FL#XF)0=?TLPCGRcHM^gaJ+3K\+^694.3HWQFT+4c^Mf>OSe37
)7@gM0(dVVF6+41^;/a,M0G<+cA((aBf^8M#<B<ZCQ?<(Z5=JM8S8aW1)KE_L1_Y
_IT4+c@>;RY.X>JT5]YfJ=^5:9fKXag6E&aV1>f.Mf(K(#V9)a2+1ccMS6DP-<_d
D>(7+9A(BGVCD/_RBT&,<9W#^-3.&_>c;Nf(@TARg9_NbJTeL0OHOU2TKfBO483X
>ePU)05B8M1Z6,3ALTQP_3>fID0)A34ebJG&Z-::3SW\?AI52;Cc:2EX?(M+8A9E
GBU9T5ba(J;>4>8#,a,QLJ.);Q0RH239@+#AME/H7LNE4[[Fc(ZA7>7G8@e^Rda-
(RVLM=0JY?WFP2c:BN&IVP3f463FGfP<20G<R5[g=@eLRIa&Ub.:MI;O<&B95FL\
)HVES#2ZceeaS[eMd0IJg=DGCRCJe3/4A\2GFDBJ#S-8e>53Z7aS,dc&DP[<&6#.
-K4-.)g1a1[U#-MGA/PeHb40]M\Z+e#12+3DI>N-C9HI3NX4JX3YHgAN2HZ2BB;3
VZ<,,YE1Z;/#VS.567;GGKYLV=aL\W5G3;U#a8IW.8dX@;PgSYN/,;R9Qc[-:8X6
+E1SY_:RfS<.QMTdF87Q\d05gK4#gDFME=HMU/Q7UW<Cd[)V<cR-EAR+<VW(4>H\
d.:0#NO6LZ,_OJ50X/EVC[#:BCET>M0MN0\&0LfRM[O#P8ZCM=M\:/\0KCYUCJA-
d.@91DG4>EI+R@a0)?bFAM;0-^X_Y<CK^A1VWC/]E,T=e&#J]^-Uf1?>Ub]S184G
F&;(&d@JFR#]WLB?+0K]V(+;<9JPO6?R_]SH?LCf(BC,N=4@Xd,5f7H0]f8276U>
6W2;D5bB(S(4S#[]SYfTg5>63:UAdR&0/V+IMZ,0KeT[&VNg:UDQV:U_b-HeIEU1
_b4I3BG3-M^+S>O;(d68fH[6U/+K.XeIKK//F8]2e9:IcL:9gKZ?f9C0g,UBUV)Y
W=9Cb;9K<GgOadE<CP/J=LOP1)<OJ1YgTHEgG9H1#JC#Y0JE5JaJ2;[NHM6VW/VY
5JC0L]dcZd8<W?<3M:9GG.#N1:eAX//OEQCX2a7UFM8IY5I3?S&18OG-X1UNM@U&
VZZ-&2Z+__>J+dLBe<_RQ;)/_@,SgJNRF0WBg_LedYW.T[<P@M\.C&?fSER@8K]-
F&BRQGd4Hfe\[U&F45NJ=UKC/bNENFXT&>=]Y=)>HO7?Y(XWG?><6<Ng>M#g4ZV&
/eeM&[g\@.,;6HAD5[1-8-eFHM..\dQGB:_NK1DRLV)ED4ABcS;X:>faFg93g2V#
;BCaV[&9DD5CPO&(W>Qa+?OW?/Oc4NF_M4)d6(X7/(B;KF^LXaOICHM1&MIKf#WY
(/TDfZ+[S19d:I8;-H,;E.Z+:a-cEQ=YK&K^C_NX4(2Y8@-(QO^/O\4.<cS/37(f
+E1?.<d32K.-FH6e:5FD\?STf_5]AHJLTIL@>G#gNBV)/#@5<N]L[43_GNSD.FXY
[WN-H2L9UR]?6)HgIOIDf#Kb5#@OR((AJc5]b^?)@0Q&-;HTf5LEU00))8=Of@A#
aH>^XaBVaD.a(bX.;e9?0S]AT@W4e/]A,Hf0D3I&J.)G^ANU2_g-S+.b0EIHGVS?
TZ5(M6N0R)<7,KOJcgL33K-C>Gc<?@[R0>P#0YNgY08SK:Z&A0)7Z=97?d#CI597
0_E3,@H)eY?9DdRf.4^[H/GW)(1]SJBMHZT9P^==_]J(aOA0/>BACc-J^d39ccR(
4?P6B7H_W-)<J3DC,K6fO;37B<,]#+#IE;HY@cQ&Y38Q3_(065Qg@/8eVJMZ#Hc3
714\2a[bS--VK:QeJG+d)bL;9e\W:K5AP9J8^_JYCV\,Da)+6-[B@2#KPF]-V^]4
:O2C\)ZE9<F.W=(ZJNOLG&23IeQ:eJ)&B5X@?)T+38&?^)]B2-6fS?aQ2?eARX/\
F)b5>IEg,3gN\C6f\0HZ2?WZZ7(;_?fK1TH=^)C<0<HcXW0LKA)6)<=PF^:fU36@
6?X9]@33P(7=DGTL07/_Q/6&Q79KdY3_a2g.WfI/4)M(cg[?U6HKB@_-2Z1c?@<Q
;OD]+f,PWe(I>J_MZ>_[(Q/GGG4eLDJ:ACb&eZZK4[Z#G5B\XZd]Q)A#?Y1Sf=ae
T(TR.[T)7EBOKHZ_1/U,f-+A>M+(VDbR.EK8/e9e_)-)bCBbA:.2+UBTaa4\F0DY
C@IXJR[G9W^J,Mf(>HHM)8J77;:;MIgd1(>HIVPKg>2aC_HCV,@I9f-1,LgZI]F8
EcISRBL8DeA-c=IPdfUAEDIL.T_a=4VT#,PU)2>K,#E)??H\G?EVbOV2eZ.eCE\\
U,8IS7<d4DPUcH6Y,LLGaV4cR4TK\Ve((IPA69T@6J\2)^0(1.SRC_DF@4ETZ6G?
(OAgfJI^:M8V6G^MUc.8<5g5ONb/<,SX@T?2P8=R[899TZ54>UZ9N[+.:4a2YBD3
JY=T&<K81:1BdS(g>dAb9Z-&f1abJ4fJHg>62Z>U)DacP^U46]^X]QXb<GZ;=J+K
YDdO]1+aE?._dS9UR_CZ_#(91(BF/WPF-#E/XXF1U98c:dLHK;b/AOE&S.b#+eYB
RVXRX)XY.<#>^_WOW2/MKFXXT)Rd^e4R.gCbfE,_J&]#SgPfI-(E=SbKUFgNSM?M
/FWNPgL5_U2ARB#O8[6D=6Q,fSJKe@#&3KafCG47;VfG9gIR?.G,D@3DQg#]981#
-5=\OJZX(Q-Z2[L15&0#OgFcJTe<U-;WXR<_T.]X(X5HVF@8\AY4S2cP,8A96OL:
V5K1[G6[Yda[U8[W27_5B2>SSJQg&JF@U9R8CcVX<0>JEMT;99U-2Fb?dK?TVK7e
5.R<IJB5/AK,<gH;5;7-5L3;O1C4X?Q7^+DOP4(3\OAHH](RFJG)Sg54((=AWd\U
g\F@gg?M-/[4[.cG^8_\\FfJ\]VL>F:=Fdgg?7)->CZ@gC<LHZ34=5)Ya[#W;(RP
?=LG#We/&=/R_]((+D<KV.<H&aM:=8a-2D>e0FZUTMA4R-K.eU>#[D\@=5</ZJ;(
&[.:9#,S66)XD@6Bb,/;HFNB9Bfd8_KCOcPa6Z70[JbX[\\R3QG0<6IDQ^gOf#K,
)SNQgHXZDH+6C-::W#S>2S63^f?H6J/868SHFS=CbaG@:1Q4N+,f^&CHE2L67Y-+
35Z=_MWUXR(NXA2IS<Obc9,-bQ(D7MdVfI1,f_E.O<K+Ef&8:\#R^2.A@Lc+7:0R
g,Y:aETCE1d,NfB6C23-dD8;L_B\bQOKHVYLFSgI\<,F&bL\B)e;X_BWK^DU:>@F
EGf&2RV(#B[XMg]f0H\e2CI,HJ5Q6-^]0e[@ZJA51P_=,G<8ONIO6IB0&3Q/2g-R
.Y;a>LY?3D0C5TCE:TbI=9-[+d.5C#9/5U)I:e],IYe)-3EUR8dO\D&f?9:_UH[1
QRJc@B;8#YTCDLK\1@U7dDPM(e0?H0&3dD>8KDT+FR:)(d=YW1NMg9-MMT4C+.K-
R94&SF,7;c?.WOc&?7_MSJgA(5)2B=GVA>IJA)4;(VI#XN(#WD=A>=U;f(J+VW:g
Q>#^<CY6P^9/1YH6X=f,.HF)[G:K2_#;cGJ68fgGg,LdfJ1FEIATO1(9=M2C;6C5
P25#RQY_EcVdYe]&+,6<;X;G8[@-R)5FWLX;DW\_1DCFKGT+\XMU&IA01<OGA5H9
&P4D)PZK-B+62F?(bPZJWPQ5TTRf>-)=Hg326MYO44gT(M.0);]+J@9SX2ZA#.N[
0UcJLT+Y)aQ2)43N69WBYBS2=)FLd>2SB\N/2eLMeb/(/c<3@P1T-VQb:EUV_bY_
.31J-;-]e6T64O>^g@e7>@3\T/^F9?VE05\PHPa\17Aac_J&T+IQ9NJc4/gW3FBg
1KgZGV+_-=\:L17S:[HUYg<-7^gL4W/GD2a&RN(\;b)-a1.2,5<YcGS8eTJ0GTOg
,=V=ZZY/OBRcd\/#UV=c>9:WEaR)GHL3HX[V;M^TU&K4Xg]C5I-0OWgW[2#=QCb)
WN2BcKU45+--T6>GH>c1]1Q<Zf[.H7YZN;PU2HYN:VL73L4M#8;=,2\=SKe5L+Q_
U<9-_XZ=\)?GT24SaB@dCQA#S(?LP.DMO?=TebSN_9\][E21/HK1<?[+T4QJ9-Y+
C^ZbMM;=RW:YA)?gB7NAN:_LMb]FL3Xd=Sb34IScbI&87U.(VaJ>Z.6?eI?MHSX2
2)P:Z.EB45&dEOHEEP^3,@e[:G,:YDGL9L9]SI^P:O:[_.HaC,P\g1TOA_B)6&P@
YH9VTe;#Ef?PaUZ_=-HVI5N)^VOJ^;UDCU.TDST@/.+7OG>+d?P.IAIFGX)^;=)J
(S&[IG_CV.06]S_;]b@+d(^]QX_NZ,)\,YSbT3#TI;f@V[dgX1bMTCK^[Ug@87<_
AW@E(8_YZJL-fBI2Ba#0X@C1B,1;Wf.GU+2K=D/ePb5B\4=-9[We6N;)F2>\b1^2
WY_#gE3TGPY:,eX0/6c086OK_;BVNV_6.A/9<@]OcERd>_@[Cec/=E\DWAL/Y)=4
Ob#7\6?@B-Rf&NSGT#\M#L-(]VXMRS(NGP,^XA1#TCV(K)K&ObGK3=3\@FD;:NgW
DGPA_(FAFb,RN,T-E&JF_YI7cTa/IA#9Q.Y[Ac/;//+&E3WM+@9)b)[)1Q)X.dV_
6UXUKR5a/cPfaU3SY;2DGIe,:T(??(R\>)K(OQ<@<+aFZ.@O;e[=?Nd<5OX7N.(I
Xe-<O_/GFRga[NRd\YRZ89.9FIMf3JDfLO+DP]?c6g716<\ULRcUO)Y++>Pb9>#a
ZgME;VG-fCPg[8fJ/40]]@g[2?;K9M=85O/YfBRXK4#=<dL(HLeM#9X>I#[?)I9\
A+W9EX&\UgCQ([72N[>\bG3M+6FUfb0RI:A2#6#TPERFOcFU]5M@KS.^2)-3RPCI
U?YMIOBY>T1#HGB\#SYCD&,3BfdFB_]f+#>14<7YHJ(RSRS<EZ(0ba8M4B?APXIO
?0ZPfG@#PO_V1M_0?[A083[a&8E[676V(AY\E^6Q.T<9T5X#4K@4\gWWd[3>RHe[
0;6^b]=77MLd\#@;3G?b-O:_cbF9\,G)ZAV+_^-G3R<Z.I7G?MX@0QM+g#[AFBEZ
e7Pd0.deK6H:<+RI,,#P+BRYDe#-Zg:T;(c@)DT&G)<FBcaSINFdA.,f-14fA)g>
@CZ863C8gE/2(2/bc[b6Q/+Pb76bOTgSe#BO48[eeS58ST(Pd)cNgCKeLT<X)Y4d
c<G0WEXPe-FFR:L&@25XeX-0IC/Eb)\XZE\HLS[S2#SY^VZ(0/D\a-I7+F40BNCW
8T;&ZcSeARMOVC\a/[6gI@GO;NLUSF83U-a0aB(XPR>Ee?W[DKBFON;PI+^dPPCb
,5,POE@7)a7/_N>:<RMX17RQS+@E4dG3,bS#_6bG-WGQgETU@];WONFWd(HG-@#M
82UZfJ3\RbLd/8_d8)f<cQD&HaS,:K7G-ZXE:/DKOV<KT2[aO+;55?/97W&5c?7A
X1(Z=AK&>(P/gJ0TTf=#DaOFbHX9\K&eR]dPgG-0Tb:XEf&4+)#bG7b1_;4E(REN
\?D,O?I588B.]U8O-M]8LgVC.bReN1&Rf]/.DB>F7\-0@/C65=D_&c])..4bBK31
]Ce\c/^Ib;IJD652:37OV#VM,:8^=#?>d45ea3cDBA_bgJ.9J.DV3:1ac9Q1G^=f
c)EFZPJYD&eb:4?A:X;_?V[7LB]2S0_f@__I<#UWK,U.cRPMNQ/O\b?L#a[X?3Rd
QSS)-/+IR/dZ]>,#-[YYJ2HbRK8W;[3F:@5)0/?I3e8(05T7DY=a<8XYAe55;X^I
6K=\&94D_Q+TdD/cNdC705d:BDQ=HDaB/;88503Y93.Ic=>L0]NS](^G<]OB<g]d
bUN)7@=9KT\U^OM&??FE,;3\EGGb5]F0\HB;S\G3cTW:\#.MMMH22;dB?N(OZ.Z8
)96:[?Y65B_O=)b3(@KTO+LWN_2Y2F(74DC&(5A4V;3b^:#7KbI;QK(97E^/[7M9
M2Ca(ARH&cV0]dSM(/gfT?d>0@D/>BHXUR?\7X^@D4UEG\@_g.PWNZK:5&=d,-ZQ
9g;.K0QNGb40dbT,T<CEcGJ3W:b#HeUG0Nd?1]5U=JIe6c3c+S5_(42G7SgcVedF
+NKVY-MS35bW\7b^Vg2/\VBC?ZT:R2e^C]e7_W3=Y9H)_G+:THa,<ZB1QPGEaE(J
GR=WI(Q6Ge&37C@[88d1JIC[59UZ<8P\g1L,<\LH4P<N6)67dE=:EON90<)bTJ8g
HZcQ_KaF:XAW1a2Jc5Y0@EWDg_>A[GM]TVd],E+bPNg/M9S13J/)4.^F?RC48f[>
^gdYJG\S;QDJLBKIdYM3+cJLd]FT#@9gPc0bS-V3&PW[R-GE+2.XG.&+BFg]Y3LQ
H11RAR&D+9ES,VUDJ]<2K7P8<#B:J1^:>0-<g>9R.C;<L^;BN/RL>>CV<ZHSX>X>
N)eE.]1W,<J0.C617S=+f\.^4GdaXKE+2B>-FA)EeT#:EfFK/:\?(4eBWB()a]MX
,_O]EQ_E[FW2JR4XY)77,aZ#8D)2#OKL<:E7T5_H/AQ?[.Z4?2H4eOd9T2/5S.G8
X6<<R1LbIJ=BRK;=UY/I9QT.1J82>G@[dM,NE=7f9aJ[[gHD@QZ<X71#d5I:06>O
HbUH7D(9=7CZdV)@b/OH1,M:Y=L[QXUJ^Z/C&a2Cf\ZaafAP,.)-[:QgJ#AGTKAd
c.7SED/bTdS@^c,52Q8FN5QST=;;/UB=dA;,(W.F4X2A8),:KB,^eGSSURKZG003
IS9,]DP8>]&KK\Mcb<d87Df\(D&[eJD<A5?cNYb7>:KDc8J/C-=,MJbR3:>C8:J)
>A.AWL.GBfP0B>X[c,)bNTMI/ES>?=gO48IVB3/&Y&);@/9L7JaOKBfeAf;/b+Fc
\HdGWc2>0b<TH[)2dMPe(A]:dKe>3HEOGF^gKK/WPa-[DX<.KHCLUcL.(Sc<HS+0
32S_0PO91AGBD&gLI@gLT&Qbe\O652?XH1=KH8SY-^aG8LSR.M_>J>0MMGFT3>:F
R34?F,+O8>.D#&&PEG)eb_fQ6APbYRAK5;b>T5J@cDbOW:9RNb-.C>BFIT-1,J>]
O?CJD>O/DX63@gbL??CWX[6-_R\2/HSW.RI\S/fY)e_KD/]FgZ8QL\[?<=@ee)cN
/WKJJC29&dH\V0Z/&aP+=H,@6\<ZGR\53LR&fE7B8(^W^T9LHK?F(\bTWf0<1@C&
KGI1cc./Af<2RPL<7HGZ:Va:^?gXe[X<7MEeNa/cHgH3C:ILgdd2D/GW#A?#HXJ5
NC-WK@cT5U<<.P.I,TJIM9Y6T>8b?aZTBYX>?S.57+5[:4S9@OM&Q1)?A/UL,Da_
.]7VaT]VGV)adOO06YCF3^KY@K;&6^-K=(XGJP/e(JaBNK=<<2\E,EE1G:BM7V)K
9VJEdbLTU<]e8M=?_L:dG8Gg^A1f^EI5(N3WAL6XOB[2g(5f:SF?6[B\bacJa1D#
ge1S4?gY#g]_5S\K(]USRL78<:TXV(AN3P@^.:,_U6?_?dC:.?-ZD]4D&6[QLKBS
;.4#1W&]7#[V.bY):K5e4>9KP59?J\.#;K=4cNV?4.=C1cI7CG[7=g.0e[4c=+6_
72:<7A3I3MY:7U7:H#RI3O-?U:^Z^W1A,DgI<].gE-=L40T]E/>R038N09c9/g;[
6XD+.^QGW0U74.a&HV]2FP]g&_=C9^.Ud4<BB:-&eFTC;V<20.8c/6-Gg8Z7&9M#
1P-&QY?41QE0FN48<:]1TZ<MS8E?.e\7K0GXM?F-&2]aA(g6O4O>[NNa#B\3ST;A
S?08X&b;HgX8&bBY<]2+VF/9TSV?5Gdc@TFD7X4/QHfFOYV6;&>0gcT98MUaGWZ9
c<5f.\1<dN.#NcP-c,4VQ5<?RFM#5SRAT031#Da<[::)RNO(U^f_CMaUW.\C#QT>
UYfIA@2dHS^\K3aG.M0#K:Tc)EFgKd2\0GJc2OP;^5X;M<OUS9O;X2ATc4)6D=#a
9[):WT#:OVEc[7S&7DI)GYPR3CUPX?M>K,a^bVbM.5SL?;5-&_OOUGJ:WTJJDQ+M
<(HU[ALdb32),2R50I-L_8<3d@5DW)4F]edR0A5T)cC=8Q->cR_V.E.D])<.@a(I
A2f,CWD4b[.?9c:?N6Ib3\Y#[NaTW+)O2,07U/gECZLORa8cS-g@&PcPE>-5GA;L
:3^)BP]N_1,SK+GEV4gXHaWMWbFW5GbA:-I?0DNf7&MHBT]@KEaP;9-F0TWFB\_(
SHOD;d(a.K<\cB8\/[20Z_3d;D6C5+7bE5Dcb44@#(ERdUW53fU#b7C3//R6aEGa
=D94?dg:DN(LEJ3R?]U,S5E#1UD)#-P0F.4=H1@eg2[WE>FZ(A/0&g.XL7O<[Gab
PGM9f@Q3=01A_AG;0E/D<)5ZBSML_>Qc(661XI.4N\^OG(:dR<R:Y^P0UP=S;(=Y
5[@2&>g02bNYS<,gFX]cEO3GPMHP+Kc8abb/@B9EE]/_=F+>dgC9X3ZKMK.Pea:J
O3f32C[9Be7]BT,M6,7g,OY#YVc>DIVH5[VI(F.g5Y6PB,391MCU6Z>&5TG)N&/N
F2fa2bZJ;<C4D@#OT/>C-KC(S^RR9E@>EU(D&9b-aTBgOO<MJ9]aE-1G<T<F+5(U
0\3L9>QSDL9;,:\U5ec,\9g>\=#Aa;^_9YE]SdPPBO82XDL#TR<@&Z);B7@QRUDA
]/_;ALMZHSN6fY6eMPY(Y8A>R+eXIF).,.9A)@g]T8S2UN7c[^bWWX;@W,(3e,Nf
+B-AgTD>NH/L&CR_@9[>5/f>56E47V0O-XF((0\e,T74Z/3K+gTWG\<W(eX.Og@)
\A;Z0H=)@6]G;YW=)Oc<GJ#6&OSf[(d+bSUfF/Nc4S[ca&>ME/gX_NS&LIQM0f9+
e76)Y&\\)SLPDNM;I8LcFG+.6Ea3,AC(:\+G+9/gCC<R0OEICVfb/=>?.CabgeLO
BCf.Q-GWb80HQ011eVN6_)eVM_e,/@(E]=M??>S,;^[3f0(/e:0-?HP-d.BaPW;R
RLG2[Z7&]8c?)L<>TXfL@[MR53fW2a>8[S/]#NB+Q@9&5>.[#7]Q>&)A.CA^8b<&
W@F:M-9&WR<[):JXP[4KZ?4@I@<)P@(e:aFEBbDBR;#<1FRS[#JZG+LE+E==6:IR
fb?N4M2FfFQI])M0O\,MGQe(\Q.<1]5,5S,;>MCV)Y463?I&N:b\:3YA9XD2VA)#
NA&K/0[^63^\PU10?A#E4:6QYZ12bU]@F[bd>G^K(2:@]Ge/_&15/b9\EQZ#KUe:
&,@^6e7H8N>LS;OWV]);3IX>GL4TZJ^VFQ8,d/1=cTA;QNGBCabCaEfgIXFTbOCg
Ee?A64OM[c&ORP?e^P58d-&aA]/@<V/5ed-J2eIPg)J5V:HXJf)WXP>B_#\66)E_
/e)33=KWL01HMU/R:#7R_:3/G->?1--?PIBbRI6.8U[/=C;UQGg;5-G@4Eb2YVWW
:R8e8M8U<\DbK/#]9YW6Rc5c+,N(]dZ\#S,=c:VUYPOg4f,AUbF:Q6EAQ?O@Pf0-
EL\&GQ1Q:RdLN#b+S]S26gLJ\3Md,QF^7P<fBg.)(MP(E-/8H<NM1SSYc>2)L,S5
NQW?JGDHf7agZA)51L<?458U<J4GSfd1C(-Tf7AEd3#SeZ]PZ,3\YDbBe7VOSVZX
eKP8D488?GN4aXSTC;J(AbZGOS+#]W\fBK<B8+_S3,ZNf.,/W\f:4>(?YLURcGUH
76#Qa,DC7M3e^VX[#B,eHQ)9YE>/g@R&bBKfaDN/3[0&I49=FT38:BcX?6GU@cUK
]ZBX^P?^(R]17V61R:EbLdX/25XZ]c]b._)OPHQ;@\Md;_4c0-Z&A/Y249/UO/[T
R:.(41N\H>UG-(@\&G^PF.[?&PU23,g-&a2K=TB]E]D7NL&D#=/gfQbgS=Z#dL#]
XD5+P_R3H<+,62).W_A5_/7P8V)S7Q:d=@+?C-D3A.,<:&I0B)MWbM8>OVM&g6Q3
]J\[G3+F6fLd1@3-0=?d^9K+&dZ9B&&6(UR>EF#fQ2R.Z+)M+J;\-cI_W.a+geV(
<P/J3X^P_+F>X_7a#e&_:XR,F_Ja^MQf9FY_CDW+/3K8f66&AE3YGXM:7T=1eQTK
UaY0BCNRE+RS2]KB+)-:)AXfb-_eQAI_5\5?d,a/-O?-T(+T9[704>=\D@W1/P24
a38V>J0X&cPfZ<V9YeVT1HJe&.a(O?CHRDML,_[?<53SH=:cRA6D_Og+CD6R2/+@
GIW(N2b9f@\4\D3&Y/SAMOd7E4]Y2\VUeTXaT+U+LP]R=H8[89\XX;D4;g@I#.>b
#0W6XWd80>\UTCOWfc>BeN15DLXb2c:X;4c;[B:A]QTV13d6F2=PIAF,aF@G#AQe
#c;0L<+&:@#R#,]O28[gA^N<C-1^@5,M6dV4^_NSJIP20?.A#^79C(.N&VD?V7-e
:gC.R3-2\SAaR<<N4\QYC-QKJWH?><:]W]#8]>=(C08>Q#ffNM8IH[8#G7)5:2>b
a4)R19Y]JG/(XFB89X89I0Xf,4g3Q,32X#M(\QIXIW[V\R;Q^BW,@ZDC\GA:dQHV
,6LN1^6f.f?<cYR#[Z::7.b3L.==+.F#59Zc_dd.0aZ\<UI0H#]P>FCIOSKT83E(
#:#0e?\X#.)J-,fg>-fKFT[6JU@LX>K[]3K>#Q1(;Cb>^gdSO[2O,0[D-,Wgfc/C
]>;4Z:a.STUKf9MPW2QMW/-5:(>FY1I2N3?MML<8?DZG-H\A<O7QX9aVc0(Ma7WG
EC3S:W&6KT4\[.b@4V_BS@PHaD-X4?71=CCH\AeO.g\8cTd2Q[GR6BGA00-L4/EY
[]egY=_S_+34,CU;RO-^G1IIV-TC]ATDI=gR:H=/\W8(d,:/1LU^/OIQFCVc.YVU
@PYQdcKD)Q+<M8Q@fFZITCMFD>F8>fFHKE85[#GL4FM84+H7L\_<#A=H7-)G@W5^
;fce(G_g#Z#)B((9[PUeXf[+9EV_UXLAZ1c#YYdAY#2V6gHW_GMf(PUS@>.W+[[B
ScP_gW;YQbVA)E(,JCFc-9NBa+HJMRIO)f(9HA7SONaUTF281)XV>g(@U-H,Eg(-
1A;]O2\fF=@YO+)NYZbSBUGM^#:5NTA)38_aP8:geBD;b-Gcb2@Sd@L(#Ec0gJ8e
J;c;IRc3QRZ5#T(b@6#BPe/;Q.D^WO(dU_;+^H3a\NCQOT05[/)33ACI(2UG14PP
&)87T\;8W7>/ag1_>5H4cc:(BV];QIKT-g8V^>E0N.>LNc#[8bfZ?=6fK1:G>A0(
2V8_^([,IF4S<U=/<Hf6fNL69B4X?75L2D=Fa5T>K.DDJV=d\HX:bPd3PH.<&,a?
aXQ8^+a5QWX;HAVdec5?2B;5ELgE#Xd[OT;eB\DcFCWY9.<1JFd2&adMLQ&Cc5\f
b^)ZJ@#&9LEL66Xd^>bB-G54LO/Ce,#A+B11YeV1X/OXcHNUE;<[e1@)#=Ra,TSX
)SD3#W.&2W_IRTHb2_Q:ON(](cD9FTWSW/L_BWIW1YJS0LGc]TG@U]02V^a(/7R(
@^U#bO/:].9X(g,NT)Q93fRE@QcBR8D>KDVg/UbB4WO3SU1d2D,Q&QL7GQ2e8K&D
W?#O#]0Jcb4WF7gX61DW,E]R^2(d502DWCTT5C8f1C<99(L_AM,N9Gd:[CY8ZY=C
\f.M06dG5Ea?Y/2I@U&3bc@g-R>V+g^U):54W:/9EM^;fRbYOA5\G\HZT6LeKL+d
cQGab2JBO]#5AQc)FZ?@H13>7;P9Kf5e(YefQ&U_[245?FFgQFRgT)5E3479N&NB
K5Qd<V&\9KA_Za;4L&J=[3d=0)EK;]H>P5.:VX3-]?cQ:N?5UMWQS9&c+(/d^40[
FGJ2MDf]B^>A\OHecL61E9L=-@g0GecaQg#JFaB5<BeV8OUW\_PJ+J9;XC?+S<WW
6:aYAX^)YX^CC,V+B<RgM)0[I17C1V=YL/3.dbF9:5YUE(IBBK>1[;0\.FDJ+-)_
89&R+aS4Cb08.f2K?dS36gDWc^gB),(#CefPDb&BM>;/[2WTO;EE[c5Rgd1@,5/D
=8?43=La/+^ZB<&MWd08dYf\Y1I6Z?U-8RWVPZ3<.S#2S2;CPHKV0Y?bf-7Q,?gd
25<<4YABF+8HFF(4O(SEbZ:@7UWf=Sb.[1[Jd>;>LTCRF>SYd8Y::c./=K2g=0-\
KYG+>.0@45aOF7F;aZ[OMRg,F4QXOeWKgDTC\/@6+e09)H7?_DVbEeNgD\fUE(DJ
<gE?NgD1)>b)d,<=J-064H^T)0;,ff),PLee8gF6CM;KUACc(SP,?7<AAL7.1g(,
XX]82R89Y-JILO/a]H\7@SC-OP<WWGA^B1.:YG.ZUe=23VZ<b(@W6:?2BQ@E&A/6
SZ/L778-Y0TMc&>-FX,TEZ;Lc9=K-^6PUS8:IZ&;Z3/E.H,I)C139Ud+GHafT(K>
Rc#\:Z6(UP>=;YFa<^ZCb@fPRU^#(gO4/QA9V<?_J-OP)]aH=UM5<Y-/E9.dZRME
<g+O7>H]37CfE9Z^)IZ4=/<55)OeMe>FgP@&X#XK3TRX&\]3L/B5bAY7.KQ>=^bB
CRf:.A/L:&4A,D1JVSPBf8@BE).4b-ABN^edECCdU2G<g&.6]d4>Q0cZb9<>R=,I
A;g>f5([/W#eUIBZOK)9dOE.dG(A1:4DP;dW7?/@2?e]5YKZ?\YEQT9BTL5R7]7I
eKEAPO<Q6++5\G0JTKNF2UEO_XL<X>=D)_b2\V;XWVe^TPS6AEL+e&N:VC[-eODb
8H5f;^=H>Z^A_DT#>3cQTU655DO)QPMPaNdBC.0C5c5@-e&CZAC\5.HK:+9Z11LO
.T&^H][,8E?dT6T(:BI/H;0M6<FA/003TRLLA2F<1f_+dC[1c:4L1V^PQ#,f,D7K
f&XF@#H[HVRR=X5F9]UV3,UO+De5\a]?)Xg9dI_+.Y8@I2Fb8]g=g^4RS5K1U?-a
d^Q7b8d4Z]=CUg\?fR6ZVgLX+RP:X;]-5+B@d?bO+0Q48]@L:DL&GGaWLaT3b_X5
SU0&D:S;DgG1S;N[LY(gRZ;a8eZSIY?N5T5BT^7]-5JeRE1R#fHeb+[WIOL@T7fY
6=)#fNSM74DMH^FE,(gP]Y:eZ?R0cE3@QSP1#fRGHaQ6]12]-MFV<U7@3ba8&c<B
^.D82a4+M:9;Ab&b^/NeZ#N/76-DXS:UGdC_8=4>(M=;7,fYWIC6&;e=QB4)GBA.
FZ>O13X(K435/RQ4&(G]OH?IW+\<>NDeXWgTbY2MR]SeFbYQ[A0a.P:6UF[X^gBP
,FNaMRHF<I;\USa,5OVK/WVNS8CO56NT;LB4>?G)9A(1V@b]ZB0]]L-Y;LIL2_gM
HEd)A0\=Lf9UXBOX_)#XD<e&F;SaXQ\ZUMY>]4#AZ;FJ\?31^a#I1Og->KZ-EcHc
C#Ug/G(FBG3]08?DR__U]Y:_XN^12<@Sg/edQ:F6,3Fd_ATdR2d#QVNPG9]_e>UU
2,)LFf:P+YM;&Z6D;^6WdT^>HGN^RL_E58.c9TFD;=:b?UB_R9/>,@ZB3[S?7:a.
)bb]_5S+YLTNf4OCHD]Ef>C:S-DJ2X4<5S@\0&-O8G-3Vb1[)Vf<b/\S12)VWdG;
eHFQb1[C#DCML8Q)X:TNQQa\e=^KQZKRWW\RJKIC/0c]cQKW&S3]2RA.d2a+,RS[
SM3L8aS_BcaKI:[\>TEOIc3M5]X)DOUN1.;<BHGN,b-02QNIf((BB&gDZQYCc4[0
7UTT7PXe=aL[(f64@&C2Ibc_GaWLV=DZFTL-T;=\YgYL_55Y+QQ]aYV/JMRc[O.[
M6^1)14g,T]aM\=;?G\XY,M<KTB\DZ33E8XE,F_ER1PL4)]VFdPGA\;R4>^4-3IH
X:A=L.^4a52E^AV0BG\;_KgfHU+SbS.]6#WWM-[+gg#2ZZFLWW/UET.IMaVO)4<&
C-4GNTb6Y0>:YeUZ>TQ^NW1DBX7=(f1UY9aQI4Y4d/cB4c6@:2FQAIY>YcbPG7D1
9Q73,CPKZFJQ[e44a&MQRRNO_f==Q@LHQ[N,Q40(=^:6f)]C.;&J/,TbS^bDS32)
L:a.g5RX&=)??C@OLgZ#27]9&ZGP=,@+4NWL\QdW[T>&cP-.ZZgSVa=ggVDO7IO9
N;JNRbLQ+MX.Da;YR(S/.Y^NO&gVa&Ta0H,bHC_&NN9KGN1&Xb3=C@7#D)[bLW]6
R7BQ@c0==\ZU8B3<.A6EP=S_BS;I0KeSVIR4](-F5D#.\43A&M-AMIe8>gEeIbcN
8AYN=</b[CP?DOgDF.#SW+7Ne0HG7?AgTId?G.L:AMefQeDYgGT436K4TD?K@^E1
J@7XGP7.F,MZ,P;DLA]-JAP5(-cVVMH3:S+H\&HOVX?:6K)O)8_S_[A2;1=<I:AS
Y<?&0:G79#aCKC_,G8=H@I#78c=A9=3@IIRa8-[eb=V2<XQJEZU>Xb]PP?T5Xg--
9@g+=ZdC9XeAPFKc5e=<4bS9GFE-V?WO7,566Z1RJWY\#_T8O3C1?2<MID_&2b(_
IW\cV+3FU:HC)E+dg]+UO_(O+A^R2VG@(D#CL,cOB5CT4Z,45-f5Cg:8g7e\CgU(
]&f6@+2XOF=()d82PJc\;5PTgTFH8S9(=0\&D#.,Z>:2F3=(>bD<a-+[Q6A#TD3P
M<D[[WK<-41=I9+:fEeVg+bagC^X<>cUJgCP^Ha5a+5[^W3-SUdX1V)9=8,eG+^]
GH:PV^2IPcbc,Fb^Kagg\0Zc)g+gGB_@gUL:2B8&E^@9H1Kg>?I;T5fZcRPYN7EW
\R,MH,Z0OeL41Y<eBbG__)[N:3019Rg^6L:d[D)5-S9]+5Y25edVC84TA;P]LQ8M
MJF@AU\0Z.P2OI6^4,MCJg7c,;&d(SJF[K:4S+N__@^Bd1HSU@K2\=C0.dPLEEC=
cdZF7gEB-N_VPZ^AdaaU7H[c1OTU=1XNUdW-ZLP)JDaU+/1TV^617N,<>T5AE<U)
R]X-]U\P0#[89<E6):/g0V(dB5]-8G//N2_B/(#fJ<\>6P557^CW:@(02c[M?J92
b6ALDIAfN=+^Q?\NR?&YQB..W4D@^4/?S_BWJC2)LW/M/&&03c:)BJ8_RN_dH.>L
0Zg8)\4Q\7HRMT-c^:QdWR2X1cU>AG96(a5P:_WKdUYT>V>&@QD16SV&/d4ZJ+\;
)+^/EWM\<#7ZHaUZHE.GMD=;-\-1QIfWTB6ZL&Q3(_c0J:XP;E;_fLKF\;OeW)=3
=2DM-fUbSRTDDG=e;eP=O?9[aF_>02BKDD.K-5\D7VZ^F\F4XS=7Q_2S9VOEYE/C
\dJ[g4Pf.1R;-9=aCM(Ec;4D#TB^(G65;QZdd(G8W+2Ta347UZ8^e(I6CC98;VV+
O##\^O=<[PE<N_IN+1>^4#:,=6(L==W8>JeIgR&R&>SG-<IH57/CW_T&7L]1a3g^
[.+>\YQS5V_(=6PVIWY8@,(ONbe4D=W>G<5<=DZ.L7ZabP8XM>80I.@9eGK<21RI
-bgJ3)U884g<0M]NBGg,JQ2K-:MH2QDX=YHMLQf71#B^GT0N#_FI5DP7O910SS[U
S&>_BU1LUgg8eEcB998SfMZ5HZ;=dfD-H=/]7X^EdAGV4P\e.#M63O<\5GL7M]Jb
FNTJ]<?SV=g7\\SCQZa[I]\,CO+\/PGP]:(<QYgO-+#[0d)@UU+c=R\,=2RHTeT/
/cEVKH)3CT8;Z2X<O^^cdJ@c6-9,\<M7#W\;-#^\,>+N,K\P4DD&UL-TQCQe^G)&
V5Mfa00#6GN)L)10d;Je[UU@F2BaeU5,F\5aY]CDB/KHdcL^S>gB/QW7@.#gD6VC
@O+]7S-O,Kf<Qd:-F<D>)GS<RI#c]877-:K=\/7)Ue1&@X#&AIX\9FKc[8:d57g1
E-JOCN@I#^bS3[XEAHHEQYI_.#YIH9U6/M41:UAD5,XCfR_9-Td2GQ&#WKe\V:]A
1HcA1BYf7+f1^a<.NbD7I[OA[&OP_LZeFdGU_IL<<YW<)S_H0B@B.RN\3L;PRA53
JSeI^(F:51POQG8J]7WgGF?;.LJQJH7N6A-./TU4AQGdeCL8?YaCW.5(H(46K_^0
29PaU?Fga[/B/_gE.cd-b(G:_aRYE,_3d.66L-KG,/AW^56QF6Tg9Q,QZD9(JYeJ
MH_=WPCCWK1X+;fE0d0d)N>F-5B0(5f3H]Ze+C+gI.,9E?U7Y5EY(?G\Q3;;X5X[
+--cJdJ?[TMB?7;K.#LgffUK:ObQ(26dVEc/;TKb1gcZ762YLNU^_L-9XfF8]B@C
:.>7=T2#.TFgSe@(<-E9)-1<;F)T)72683&#f/Z9)CN.7<V0T;J3QgcH=Ud(8@gN
WQM)B)QMc+B@DA9OS[aB&)^aJ4F5K#)&\JFHCWN:5176[)Q-;f.\3[0GXg^1)d-A
T8)_+YN#D.L^1S5,J:a3](=VQXB[(Wb5;/)TO#F?b>IV+cPH5Bf:6[gNKbb6BSFg
NFDP[Wg^,J;(TNaa:Q8SZ(LS)0f3A)X,]9bDKP.6HV.VG]82(.UTgb5a^BP.:0;K
T<OUZB@SWU2&WRN52&\Q@f58B1T0E><c-eVR]5F=bC^?cWMIS,&/>7dbTX[LJKL4
I=>E\QEPaLQf/^+>Ed18?U^<F(IF:Z.V6-?9W5.IY)9HCIX/TDTELY)GH=4MG(;]
dJ<GDH.QLDP#_(S/IT>=+7CQaN1IZGW.H_F0\B[,/cUCQOgG=[PYD+?Ad>HK7.Nf
ONZQOX>aMGS[9J=_f>20G56YT)F?YXJ7H#X@6/:^c4L3PM?c8:<#E)[W3db^;J>a
RXS>?+d@.fU.HG\&gb5d5]b-aMd.E:c.P96O/H,eb?<-bf4KSZ:X#1VPG-bT7UDP
W2X:,.AIT<-@EX]cEYD@<]AF+>:7JP0P/K)dH3H+H?5<]FCW=NED;S5A<QBffZ&,
f;35VAJSN/<+X]ZLJ.1TA:136ec&O735(Q87?/.IGPR?N)0+eD;gW9L4?<0\]8HB
_(MC4f(3#V#Ca+OcTYS,b4d+<5;74P>IS=WHgY9A/;3[TVHQ7)BL?4/;eX]9R4R[
FL::D&D#@YT;UDE;4d7Q+-bH=,[M(Mec@9Y)FK19a2.C][a:KXV[aa&9QBa4)7ZQ
S4g_U47dR.6g\bIYgB4K#UJ0?G31S^;PgNP5S.<[IN(GUUgcIGK?Ide8#]K:06H;
F/BCEZ-5^,9XMS0G&A1]^c2T+22@7c?3+fYe[FeVb^(9>O5_P5;YRCLSC3^.[a)U
G.W(<IMO\JBc1IM)H](S=-#Y^KF3;FfZME)>1g8f5C;N42>ZcSB6Cd]MFT):8_1)
C-bC_J3b.J>/<-cNX5IcGXQ4(dI=d6DdN:ESZBCLDEe))7@^:#>c#K+GN>B7L#?]
E.QCB9/W7?@b8#7XOH^76B4MI0EGHM+7<?^DI4<)?><7[IVf,bbDPPZDX1.#P<e4
RUU[(Gd,)9-J0S#Q^PG0]IHdM3RZ,<#ZK\f84&>9V@>[?,SZ+(L_K[?5M6#]VE@4
UKGS)[,=6d]774:Wb]H.>_B7deC[PRY,eUIQ_XW-0#=005WPaPeDE>=[4=[0CPJ=
X9^&SQ#O8Y[g&.:EAXZ)&I3NRINaKU&]R32BSYd7WVE,QJ@@<1SZ7HL)24D?=@B2
AQ-AgR4=g>>B.2^S?:8)QUZ0,NCSW><7dF[dZ<GM-AcCd[1YN.F<JgI<X3H4a^LJ
#:9(&U&/?cg^QdPW#(C+I#6CfZa^agLB8LIKR?D,+6VSZE,Q<d:0H[/BB(Z+1c\2
\e.UWQDENfMa]2B+X[PO\9BI<gY4\]=bI@1;e-<@PgeTZMC7BFd.?[7CL#&@>bWT
&g3Q61QSM/FE:XA[dOPV_Y@VUdY^32N80Y-6O6][KcIJEMF;[fMDGN?O-]+IOOb7
RdL-V?Q41&5DC]-_91N]bO#0dWK2]#?AaL0_.JF<I3COC5d2+f=)WD;=UA.6CAM?
6,(CbF7+O[5_6#A>Y9I2-HeKeR1a4:dbC?d=5U>N54,J6(E]>#G7TO1e-[KLf]&1
9[9c+1?c\R3:MdZc/\N.fVV9J&)<<=MV].=0RO,G3ddFL8;Y;?XZ,C2I^cae<AT(
01E1^&+9c/EbZ//1Y<1DAJ>31&7bQ]4PEZGO>6DdbdG_L;+Qe+\/Nf_;4-&/FV@d
O:F1I9PM+O<AO23BO<461HFA;R/:YdK[Z90PN<&Y5[_=#FG2+C(-PX)CL3\@H-&Q
SK5]Hc)I[KYe\c=JBJ?A2,EA=NaEgU(H;W[<M/WPXg@DUQ.3Ve6>g<M8PNA3JT&^
N)J0U#V#PW[T,e[/G<0HcUDYRP][X,]/fR79RMNEe\/HA9.S(N^YU62=\UW&EKD&
3U]>d616LRW2dNP&7=(ACbD1?U8F<RUBGB^(R6X@S8e=&WCb\c+6/d4#20UXTc\a
F<;]893.N#fY+OL\;L#-YL.;/H2V&XJ<=B43,)U<0N<&Y]4,T3/S&Ccg_?@O;+&c
M(Kf_8-_Q;#;((1d9TY[+_I_TO,b;:1SfML^QL(eSBIK137,6#f#cYRCg/Ea?#X/
\Q1#Y_DJ3.?(QcMgZ[#><K\f;UI)Ngb3ULWQ6+L1^EA883FMAML(JBdWFB1+W]O4
E/P+0M[&Wb3B.d1C0D<-.G2;88;Q^M9RX,[;;1K7PGT^IH,J<.OgQXa<+,TD^4DS
(N7LYIgDQSb,>TM6P16,bgJ8F6f?[=2,>\O.A/O;^Q#:N:0(dT:PX2]Z_4C03Ug=
dT.DZ>O>A)KLZfHT(VOg#:1fV:Mb.Db8#WP-72H4X<M[-f1YR5OU;H7V-9B;J3?3
<+3_W@/2Z&QS:1d4>\IaA,M9@+_/J7E58XQ3b#<7=++K]<7Kc5\78OQ=bZ&(X/]^
0<]FOZ=X,@/&6[eK]@P)4bR,<&)5B>P?K4A+cY40FC4_aT/7L>K^KY31>D\]^0cc
.S8V+HF71?>^1a9cM>E>RO_TZM(^Z2+>FQ>(KTVX:Kf(+X#I6MMB2Q1RJfc?0?L@
P]S(J3/II27556NKXCeV5^.G[WSW/B8fI+bP6+@KUO2ggCKcddK9PFZRR&<;9)>e
_g97:4QI)N4:_S.6)DM#EQH8>K6GCM2PNN=4N:ScaW)]d9M;[9.B^B&MKWR0NHO_
UR+f(XYdIdg6/[e=.@+N<]TRQ])7<NcMXW5XOI0MR;JfF)-9ICbQ#I6NSOYWG<ZE
(YHX?a=\fb[=2CNAJ/4T70=.O=^/V2EZ\D-QdM+WLF\g3^aN.9b9/(A).[\(g9IE
LK)O8+gQVc;b9M[J?:D<W>fb/.NAO).Jd:dDD7D0/3>8M5;]&6[5NDBD=4W(BMga
HBMTV9D3c\L2aQ46KLCG;ba]RFL:499,,<UJ[;/6=EPX0L@1R)0<#bB_=Z>3ACgF
2Z7eJa#Z4:UUOKQ]+/1]]^L8RT]WG6H7FC+WQT4M_V]&VJ6YL-T]-)Ve3f61FYZa
=3f(W+e[^2DR.^=eXQ#bXI<9g+,O;=c_D@O\_A;)TF]=U<;a6>=aX_@DeSR0^)]S
MEC:(#gP9X^-]J46+;XG1X+5\Gfc;Re6.9#KX?4U<)[(VRf,;31^cc\15N(YJfGU
>_2UN)74;fE.Q-&99WO&5]Z@OQM^gTd\S;ZM@4=d#>#V;256EAfZA7^8<5M1SLC+
XMS?-)?W(0>[_I1B7&W+L6M/)eHB&dC-L=gX9CbKZX4OR^D\RSFg#&;<a<;Za>1K
:-X#3bf-]7=Uf^1E6U;CTBdD.A8D;KWIR@B>:af3B-P<O\H6WegXK1._bG8d)_X8
d(B8)6E?5FXVZ@WAYYG)I(BU;+/KC=D[U4A]Q07>KLC5cLXP3<>PXEQ0J#^Z8\cL
#EW9^7,W/f1MZW&LN\NRc4WLd-14:eWWX[BSU;6JU[-#^0]3C5QcWHEVN#S0eWD;
#:T/cVL9EO65;35M,MNYEe#+7)5/DE0B@M)&d?5/0@:]TD+W[dc_Q/OZL7@@R.LT
9\N/:J(TKWS2:LUROP\7Q0=W?J6UH]G4[Mc>F3,+f]&9eY[^g8#UF?Tb;cL&+GRY
4,WD7>@KTaNb[Q=+36T+b[d-#I>YJZTR(O7<0_bYZ@OU)P2^Nag./+Y7aPdRZcR1
a;cWMG5_#).f2-NG:[&M]>V,:5bDeAESWC^bL4P_V.XM>GDD2FP@6)ebId>LTY3=
+<:e0H^Y4EV<,5ZWFeUJd2+fGC[@]H;5),>T](YXeWA6,DaDF325P6F1Y:7R7Yd8
=P+\0OJ2(1OE,dF\+f?^P_]?H:[HLcgAS/]gAG(X2g+fK.cU+\QVV]a2)AB<2Qc^
;?IU>S^R2Z\^])_Fc(S:bdG9ca605Q^0#3;QX+0bRdMK0G3SM:0<a)]94&3>/B=9
cSX.SI0<X[YUD\A@eK9JO=GY7@JSNc08/fBE-gb^47IYFP6XPJGWN-Z@&_cLVK3K
&:]7<2?>\-NL^&]M()6_;2^YIKYNg8R?2F6bJ1Gd=8B3.G&:6KHbEG==SLG#DE6S
dJBa?L8QddM(cO&VdS#SC=RcEL5G@Z.J3?#Hc.VO;@+HOdZCaaOCTSS\&4Y2_fZ/
32EQFM8Y62LQY=5C8:Za<.b#eeI_MdSAA8>f>L-Je#Nb-LIe;1S8LL.I0AL[QODe
W5#?O+@Y8VAS[YaW;9I>28?QP7K\C4fW&N8^(S.]L]<P3>5YNUB-?4/^Zg1F/E=a
7]@0fV.20.-^BeE1E-BB?^YcRHf)_ZV;fdVUPX3J[BZZ<1V6+4&F8/8Y3XdTY?36
,EHP=7RD7^J7P-T:,bVg1(Ya,JNST0eWSO@Cd)J8,H^.aZN6(?&_T=-9K=MDFA?A
#(gPg+72DbKW,4+/#a?I9)1d2,fE9[aeQ>d64I615c^]aEJKD07b3LN4-^Pd^R\?
C(YO3+0LC:_54W4Yc(&a8WQ-V^LF:8)BPdMPLZb+I70M)aDAXC5XD5JA3K#O^fXC
1<=/=bN:eKOc\AKF:MB10:^/1gD[geMT:ggZ4NKJ7Y\1a.FRYc_X5MaQ&#Q/<O[1
8SEUSB3]f=D?G132g9Fg&G;9>eLW_J9,VE#SEcM^3#Y1g.41^QdBZHP\5f8310,Z
2&)dOC&WOYg?f14A88KXEIK2OJeOGN:UX@&HV3ENYfg1(b;)>/>fPbM@ec8)JKRB
.;K)<Q=^7J+9BHEUQP\=#YQ;^D,9Yag.^9QI=8G>Xg1+b81/ZbNHD.SZfR=L].IS
f+8?LgOI&dF4<#>KQI+&6S4L1R9;IdSdf736/XG]e.b1^;TPF/Kf=43NKN^;\1@=
A?R,]\)H-QeI3#(JO#<cAS5J.c>P5:>dPT?Zf/H=\L5):GGYZ,+V26XVDSR;96#b
;IU&DNVR&W#^,8=3d5aZ,;:O9EP(D>K=/#S/N0Z<YU].ALM:WQ<I2^DdI)(/-^>.
-#^I5TLLRY\N+\f30516P4DP^,1@:XaZ4cO\eAN&O1)JaBd#-YJ3J>=Se4-@b/BR
?c7@>2b2)AE(MgKaB5VRTC_<)gYN#&YTW]XL:(,1/<a1[&;]f_/KG5eCY[&(^4,9
[_I8dc;[RT<:_C#]V39gL#cLSPLSO3W.=[Y;\#FJ421Y0RQ4J#@\:[+1X>9c&R3?
:NJeaHSN/)4(SO&)#b19PLJ#GB?BC06LVJg0&W_D(ITUW4]GE\0#BROW7:@aEZ6B
g3+DP1aO03D\+#\[TUM&f:+d.gYR:&D9F_b1BQ=7b]G3PG5\96Lf6aV(/_9g#=X<
e<a\H:Y=1S_VX54\MROcA=N??PdER_D6@LH782]T-J)1XX\_g:5-1\/?T><3AGCa
P(JaUc14;;0J:BV6GE695U9HTFfJaN9\^7F1(+#0#G/Q-.>02\BZ/BXgD83IeMe2
2:#b5D[X;NA8:\fE1\SaNI1?XFLcQ1@3+G3;=&=+IeTLb&W?/5g]F699Ma0IcPGQ
^Y)I0=_?K090b(Xf)T3>0Bf[<O+1/B?SI?CKD/Ug?O/HOTRCZNC7]@=^:UU,Y07Q
[:VPH464aDN,3#\f=[:)UNWUg/Kb@6YcbeTEeS)&=H+,,G0YGX_/I>9]@db?+0;M
I7:C9-KC#4\H]B#5#)/fB)b)C^F[MV9>?<>Y2+fB[MC8YR-#P@7L6KQ3GJ3e[:>_
@/E7@JTWd6f\X^_dCY7SVZ2UQ#^&df9d<JZf:g;CIOKfC:2S^U=G+PPB#8dLNU)A
<P_b5b-=GegfX;VMHH,IXUfSGJ^(,R3B#NgM.E+45fWG[XY31@=&b;2WW:+)@_.&
fJf_/R6[gCe5EV.cM/LHa-a0].DOM&6@M/M[E03H+aGgY#FB>_T7gLg(5?T&EfD)
+RHJdA_9?8f:&1SaVT49[6D#:=A5f1<RNEZ]M:c/SMKE9BaKJ\4g[>1KPREAB@MO
fY3@aN3-\PcA@+_&F05@fPKE2Y.WR=ZcW)U1FH+gAMd)PA)@M4a1>:Qb(<4=?I3B
9,1/X;6GT@9-YWVe_PgQ;-AA16;SYY[dO#KCVX9PLb8BC5\VABGNP+?-Bd=?PS:E
ZH)Fg\:5aA1T8^M[1G66+KA&>C19/FMZ?DR#EDfcN7@J7QY8^,>0]Z>HSN6&aH[C
V0bZ(CbdfK0/)aW2K]BRPW[Q..2DHd@J1f1APNRE]YC4ARW][3RPMS#.9@(3HN8B
7UIA_+103(<^(f[W@PYf&+[E<LK:=(/6GRb7/gL#C7eE-3Xde(B0W@>Y]&8<VU,B
Xc2[XM&A]eSH\,L]c7O=ALI[6JHT)055>g;.4/dFd7XUa.43M1&T06(1A:0=QUCc
Y2(XFWZ2MOAg01>6]3c7_8.18VHDZPSB.8Qa6Od@Ec)XgKZd&dJ@F>XAeKN,3&gT
BW<\U:]5D6<23WQe877HWB(D8-M<GZTKb+Q6Z,51Ub^GNVTT-V&O9X_1D:&1c(LH
#PGB:EFV58M1JTbQbF1(?VMUC>&d0?&D-M&0e+H?LZAKA]Xg5CJ>,7PN&G&BUO3O
X+7(J+?TC7L4R5bScEe_6O/?b2dYY4O^d8O1UXeEQXNX#0C6(<Ugg3[&d/;-]DK8
dW.DABbZ&X8_NBCN\)74E#JF]:W(]KGOF=bWP<J>8#)V6O6-W,fS;N[b[]D)D?#M
D>P^N5[,<^G30SW7f@<1EcA\-U^a15JGGZN<=HYGR>aX49],(B_)5]KK.5?TGg_e
6BO(W)Hc?<0/H+1@16LO_ea1Y&^/14ESL/KILCE&Q_I+;WL#NENAT&TVbE:,DPO]
,+4^TeBD//W.K_@=5HOF.E0KGCH6_^E01+#+NX50[\1P@O2g-955##7ATGI]QDJd
#MH^)NJGcbKP)a2V&T:#0Y--FHS6;F=XSKFO4]US6S-e^Y.1@\IP?Gb]W33A)AAX
D;a4S9,)3GDS_:\2H7];eWb_&5ZNLC(Y^]4N=e?gAF/WaMUUc&UP88a,]=Y>]AWd
,9Ae?,^N?C>?H)1O,\8)0e1cT2(5-#ZgZ<B<99F10H)e56f]XQS]AY-cLPVVCb7A
P@e?FM&P6L.>beY)P^/;WMEaI:W[gCI2ZIH,4f?&(5d\QX),f0MSX(dB,T]NX_KZ
T_MG@^V@(c0a,1^8&Y#bX#8_LMP_\^5N3,DDJ-+3R&g+JF:f.43O8@7e[Xc&VdUH
WW+F=TOfAHbKW7_,F>MeL,B_+K_6K_g)DD;/_:dIRJN9-Z.X]V8ABDZ@I+&=V&W2
&+PVA.T2\A2L\P.-bZE<4]9d7Q;Rd;)MISTaKBSPE35@(;Y>C2)9PX/&3]WW#M/f
8I0]MP]_-dMQU9MV&I&?Q_HOK),?(AS)>S+?_ETLMXGZ#X8KO0#+O>cS@e7)b-Z_
UM(=B).(1T]B,#):=dV25Vc2C86<L&V]&L,3.#??7dZ?@4T,JKe45#K#_+++,I[R
/J=Ze[b#a)K;Lae=WUb:2KW?X&J(-ca>A[.B_E<LHIX/FNZJPZP9)Fd),E^,f60Z
6GFaX=WZcV.U&]4G=)E73GQ]a3^#gM)>bge033F&8S+B_Y1I)0U\AN2CA:c,DJI5
<67SeA/g<3MdBGC5QCe]#6QgdcPU8e]<aTJWTLda(;6M^&V2EL+g2K_L1=N1[,]I
gRUR#?_IBPQg3(c#JB^.)=U\B;/DCR41_I,g/RbfAJV?[L-&3DNA-X@cEe^;e\T7
_JK5#K6&Y95Jd5FY:.J0@M,QfKR/MGg/B0N#0?PaVABN#WaMM=bT#Q9KEgC1R_;[
eV2M4DD&0I)GHbc5_,,@FCDHEN9?NO=1HZ^Y_PRV]K#K7;C43,1.KKg[&L<O;^Q/
I:MP9JcK0SG(X=@]\7[5;fTDXfgDS,^KCU7>:,e))^-T6L6,)??R=I6[RHYTU3@e
<6;ECSB\HHWeB1F\IAR\:][cD8MgB_.Zf3R:1HNOR::#V0e5]_L2=CC+8ONe,PTJ
)_bW@G09&H54Ub2.W5&9Z@#IUOMbMd594@P6MTc-)eR1RBD>#,)OX8OPVHM>+NR]
=M(?A/+</8E@L[4274H)FF[HC/DRf71I/eX:[c?2HEX\4GG[9G?LDbNST?J5J4]E
97CFN[JJDU2dHV19/SFNcHbW)9\SbGLfTP&F](b(-&\L]N493@7F),PV>fW7V^DJ
]F?CCcTbB3PbE@EPdON?59,H[,]87;MZ1a:K21=KJ)C089_/&a0@PN?_5CgM:V.X
aV47_KDY@MgBf/#14;XE8g4H9KRQXYKPHN-+DUXf4&5272cZ/-b(4J7YTB7K-gAN
A5cQYT.0e\N>9IU\H:<(SO#YBf,CN+a(e#6E-RIORHPC@4cX8aHa#4P_d#9Kd[UD
4ace(Z7L)5&R2]5c2PN9]UI4>?(H37HF7]c7G0XEVGef&;B/B>_a2QHEUH],,0;9
=U8BQ4::6L&(6DEIg:>&-.1.B-;EU_O>XF:R1O2IU@9KeVH2<bTF^f]H^B^<6U0,
<f]=T-U^[MUSJ[H-<96bE/>>FS&)^P5[cB\FOVKLf,N0Z@(L464F<DZ<)e=GbX9f
/Q;G&CC(-X;GU3@U_J6\K\XW10?[-5d)D_?cSd_)7#RS4(gSB_1]gfTT2FeU)265
R^P-4EYfI93P^24W/8E6I5J.4AI_bBb)1&:I[/P?T^2;VA1@CX1^3GL?>O],#D]=
A/+IJB>COZH#T:X\)3^#f[\FF:a&N@g8ebDTR6)#bG<La>LP[L53f#PC/C]IC-[D
,A#=>/9e;:NBgc0QCH/-N_LSMXG@0ZWO^D9?SEE6cb&<KW)MTSbL7d3RP<+IBaG_
&+)TU4UQJNB4M(RYbACe(\ZDG]?CD=A10@A4M-8Q?&72PIS2QCO=>ff>d:Z</@&f
,IH]Q45V-3232)3TaE@f^FSYHg?.>deQG7LPf)BPM1+LC/.\8_]+UG],3d:(VTG9
4](E^&A5R.L@@@E74cY0:,9C2=DY0MN-@LD[^K_>@\I1@GHLTI24W+=7fSX<JD#T
]Hb(>?gY^M_BIBH;--GB&GQ4Kd_ZX@V\U6;Q=f3b9=>.?f5V[YPKB5ZJ&b:+B/(E
93)-G9eTP1CG6</6(HXK5&FF&HUFE=P?8R1/Ie4SY))D:)L<d2M#MFOR.[L7?T^f
+@gG5d^7M/\MB8C/c9H2b-edQ;NPA60RTANO=<][2(W#,69(feEd:J?S.[R:-HPJ
eD76[-4fe9=JZ+O(FA30B#aVHXXBK/#&1;R4T9D736VdEG6Wg96-dBDNAEDCd15\
T,0A^]&RYW.&e1MU4PG;,T_g@Se&GM0/2/fAYU0Ga#\I6LG++J\0^<9_/34=YPSH
2/_[EfSOG@4>?FgMaea=4W4dZ;&JZK]1_KKJL9b8+SbY-)F@(UW?1PLOID)NA17-
RWF?cKRDPQb1=,@[Z8P0-(1/^b3?Hbb1FdM\R<-ZJ=,X58<L1age=->&7PLd@M?F
=0\LNf.4U_8,NK/D+T3:5F3OA\L/_(NYH;gTUOQ=?(OWN?-cL1JO@>(J8[Z1.A5[
K?V?48[I=P3:d;B7JM&RQ7SQILWGP]fYd(U38Yd=XS:;J8^?X+^f/IcB>:GXW-fR
P6V.A\3e42d>BdaC,6)L^U2f/?gA^83EP@WP3IY&DUgT\(AH9a#XgMP5+H,&HWGA
R.-8I>^77EGP1A2]OOa/(Y[b6fG+)/-(B4C15cXH>_8SIBKg95/X+\)8P83)PSYf
#=:+8;9:@I/S>5OGJDCd=-F.)PSQ_N#Od4:>7fM8UZ6^3,\KOYe9UVK>e1^E6YQ?
bVX&8\&]POY(<PUC5L=R,AD.<P@&_GD_1HRB)9UaP&:d2@[66()Q?2#fHa),FX6.
f)HKE2W)#7PO=_.@.H&=HB4e,],Df/IPI^,2geQgdR?PN8;@4-I@TM7<d(+#88Ff
U=6<faf/+Q4A+:JS1b6f)JHf)D+W9A7@SSb.b-[a/R5S#LID6[(08X,BeN52gHN4
D-QZJ8a:^V,C99aN>HZ39\M;c?0>B(A1T:P4R79gPef7f(7.TDJeIR05VaC>XJGA
#,-)W\+.F^5fNQ9\N;WdT8H).VPI;Z#9PVT>OD(7WEE1eS?TL[N>M?J,U(#,.eWQ
[f3D]-V(5]T)Pf\HE&;3-cCa9d_30^F[4@2f/HUVO)=N]_WQM/Q<fO7g:ST=aQ8.
)6#5a]9B14,JXeC04JK>.6<&<XS^<07C]R1#?R5=aT=;C-e:]DdcU0G;:a,H[46J
2Ncg)SVA8B9>G26g/;=\N#=b4I(0A+7JZAdTG;ADB_^]-/2=-&UAN5&5Q&MHGW=R
5\U^<#2/?R+<DV/+=NcLa@AMU[RR4<S,>U#=8SI>MD00#4M<IS0[c=^,2\SGR)Gb
LPTY)X8\IfS^.-WAW&>7CDMCT7CZ#;&3HX3VMNYXBU2a+ec940Id4OcK;#\_f:ON
WU2[+e\0I&d?gIF3EHPW8f1.>+N1c:O_JcE@C)#/6d-2[Q6dO\]:OGdf?aVT^VB7
649eC5@,_/@\aI6#I\/g9?U1dFU;:+GZ[C#<9RSYS5M[PS^g5]J#X4?+d=Ic4D/Q
^E_bX31[OIOGKTcKB3BL>I1=.e9U@K8FDL,L#_?,>U0<GV\c(N;OMHZ85^).3I^e
0VM7b.cCLIC#;.U3TR&T0.C)OM]0>LKLP4\N5E_S;]U6^]YZF\BYgG@/Q_A@(QUX
4WW_KNf?=PJMeP;STbS;TS^M_O9d7.bA2+7F[?2,+3;88fHR;PDT3M&\7QN1RXI&
5JZOP(+&9FPdC[&))C.&UPC+]Q2&KGfDM[)Td9\P8GXK,/W3NaZDJa6G[^3^ggS?
&;?HLAX)R7C^DTEUQ1aMKb(>aJPM5We\^,HDO_a.AR,EE-,,/9b?F^CBDXL(7K(@
VDF4XK(9G.eF)N??G]3b^?XG&F-c66(,I2/Z3d?)FdG[Y>b=9DCUMC[J3=R.NI9Q
2J:(2;@AfOGZ.X-P=)b(3_#T(?f(-/D1?XJ?3Ub=&0ME9f\,F&TBJT_dOVU50X(d
D2:N45Mf7/HdHAW.6@VGeYa]bfdEg0UbR;XYA54X0C<[PcR)<==XEHV/3::-^bbL
1#c-ML0eIWgXg_0a\5LIa=[N1/(LT&D-B[@EN(2,OW]+\ca7G=89,ZZaHG/5;&=E
g.>dMQ&BHg<XUe8)8F@b#Og031BAKf=TO8Y32gB(D(Ae&NGAb1074VFNZ?H^9VWI
\.Q#bR0##:_BNJW[98Bc,.EeM4ZKAY8&Ig8RB_5Mc961A+SZO.ee74,0U^e9=LA)
[TVY4Jg:9/gMHRbIS;R#c_D[I[4De^^J7M-VRE)364GMWOD8CO+?6,Fb>B?O/30Y
fJ4PX53UFSI<3(Nc,AVSCd6Q@CO1Y&KHDdNcES,9;R,U<Q8L/^B@8-dZF,9DUcM4
^g))LJN@.QPKCD&>W&dC3\),@7<6:2W15,F^/g_),ARSgaZ+4I^>NA[N5VN._:5b
J8L[S+7H+A):#KU#Lf[b+-J7I9M/RA)X&#9?)#YX_QN(d:ZNdLEaLHa\GYc<\gdR
JMM1:R4N[E\W>a?8GN4JT2AegefM<G.\9Ud<eL#RPZG@?^dY_XNB&93DV0F;IYQ3
=Q=WcXSPN(BfB9LCf\^?HR#3R[E]RU)QK]QSg^#BNL@D7QMgLYWIL[HC(aVU?Uc5
Z4YWbEOW&(;IGc:G1U+2Wa@&G/F_OHc^1:)82[>(5Q+@[4a?8ORK\HC,cJ6L]TPY
:.@4bE/-EH<?KEA&bQ\J[SISOZLTb;a=::_S4;,;CN&Z\eFAGO?QAEE;8-5AMM1a
J-B;;_e&Mff:gD9DXO;;C4;U0,Pf>NF+^PKE]]#EcW,3]3b.EFIMgLD[dgg^8fU#
2QMH6QE3bTGY17AA3[-+C27N<8bXME++>f4MLge08aSSF(OJe79=,(QeZ7__EAL,
Rb^&?2E-)T9Q40<M.4a#Pf/+/0gfN;^HDXOR=T<Xaa/@TG)?,V@Pd./F<4QJ[(0/
^1-_RK?WP@\DW6QLL5S3WcY+f33)c3?c:MR[)db7.MW8#\&U&g:P95S5/3WH-&0;
0AbBD=/]c]bBf5H<.5+HPbS-)[1EXLTMUW(Ug2,JJPZAa;S^?64PXX0.:3cI6>Td
Y.d1\Y2S5W&+gH+IO9O07Q-<cU96aR+6?H?P2_80UMO#OF3-WUH^EA5Jb=H10S(6
I0GA99VR]#fB;T=\[OS.eU4Q,@,O^>(#MCJ57XML6aP7ZZNX7DMK5F<9V>38>Z5=
cII#ATIS2&Zeb^>>D1LVV,GMc:_.+:9/37Xf;><QEeS@I+T7,1A.fN6/B;E\L4)1
FC@KBY9.\B>U&)>8Z@@)4;NO/Na:K,d=,<HW6LbKY357LHAP0,4+G-GdZR,)>>^g
&\BQ7=We;VN)[J/SCL2\&GM-=5ISd_X5Q]>b\#N@27HE485P.H7KZeM9Q7:Z4,LP
aC1e4F]+(JCcJ0a8QT/)3I0deUXL2766TR^2,@SCZJ>(HN/=535,[(+83ZJ3;]E9
)^.3J]U<ef8WeO\2/&263K^V/Ab.-aPKB69785DYHbQG5V8?Od6K9)\:17Ag5I]I
LA3YJH(7DbNc96>KU1UMP#ff0E28-23]L6__^ReXQ)-fPGdQ[.F_0EC7AN\:@&N_
WO/aT8(UP([OH7N:_;Q-9]dTa[c#Rf\bb^)2K0_9V2^5V/U1[7g62^6.Y&TD?W5E
]&^DXdc)0(aQF9H0.CX@8?ODa4X.F>aHB6.9\Y3>8:]eT\]V/2A.:__JF4XO.:G?
]V\#cFgB)_f]@g:)O4&^1Ld0S&,]<Pcb#R,FLE+&>PO_)J3aD)#OYFb]c[YQf9ZX
IM41;7FR+]2)S,G1T^4S#78,@4G:3;D9TfUSg/+Z9-JA2X4R4DU]RU;MJZE.HE0#
>UA0/aJfLL1Z405EO\#f]N_8S@PLE]K0&5Y_LWS8:NV&1X:.WX/K56Cc,^JSH+&E
L0+U.<87OFgG6ZG(:/YaXZ&-C-[][Q<.\.4S(,60&)-cWFTebPAS;cG>d?eR7+2L
@[&/Q<e?5[><d>@VIQ&f/8I^KPcX0G1g5,U]B+F/FY5)NVL:^/\M/.g@H.cJRXI8
QOG6Z]Se6J0G?W8I4BKAeDP<VWHXV-WWRD5)<SK3c9W[dX/2B.,X#?YV/1K[@C8L
YA0^[b;=L)2I[;2f,U,VdE>7g\IRG@GJ@5MZ&-O=.Wg;+F5=FZ5Q0^Mea?\]=#RR
\PdUH7EZLbKLE-Y;/EOG@4[b47J;D?d&Ba+.ENZIEO>GX2[(Jf8C.9Sa^)F[;XM-
-:>,^Q4LL:^@25_S56eZC^16(=X.)=^J/7;E/E^FZ@F6HRCG-@2KCS/@&#T;AI^J
I9NLPZ^9R&ZNdFH8BM7XZO_BQ)Q+4DIDUVY.J]DE@YAKHV;)9L&&#L:H@L:g]A-T
6^#Nc6L<2UY]Q.27PUY6bDR#1=(&ae[Z9XM0T>WW;2.7#Od+-MN:(Ba^HCI(Nd^3
[_Z2J,+bZeb>G32)1bJ39D75G#Y;Y6V;YU^#<RE15IH7K:Q1UN?/)TeZSc&P523H
B@1C5?-E.Hb2CS9H4g)_3(gK[cFB&PQ98([GPQSX(&:@H+3DPX(ObFXgM;Z^Cfb&
+8#O\W/9Z=;7T^T>/AIP3WFXg7f7R9/KR+Nca+gH3:<U#6Gb+0:+d3VTWG:411G>
4:C7g,b.R@cP4;&Y@+=CANHb/HUL0?LYOM14C/b@SUFF2=CBW\f+,Y+B8Z>A98Wf
eQSdbD,-?N:\WP]+>;KN;29:_Z=(T4_&4T6J/f#BaFV2X,0[5-aD^P9bY(6ZBH)+
W\_:.Wc3dA,Q.WET4CA]Y:WH;?S::A??MP4(,aADb.D+_#c+^>cg9VCR3+<Z#d?e
+J2<SBFc<3+5<3afTP_UIaVR/_?,/-b7<OGIORfL.[T\^V/Ce8)e\6SP[(S386)+
V(7G[aW0afGSU.=QTa6=)D-CN-TJVT4c]7K#=DfYb;N?GXMYD)5D?URSf>V?5QZ&
>a(L/D08NT;59;P#;E/Me8-&fR]5(S)(X=/F)@#<E/@b3Z4>UQ:VPC)gH^4S1SER
V&8B5^cF<,)?&+f?,;e3V3cU4T-L-L>64Qd#&OOR;b:cbUSFJLKCZA:bS]a4/=J6
4>DQ<?QV#<c+FCabR5Abb;CHX;MQAQef3O22+(-D./4#O9eE<R/A<NPJeGVf7LJ9
.ZS4;VR[708XR)-?KH+Z&C7fB1HgPG:@-\3a,c9.(II+YII2A7eff&>f;I_;3.,3
Ia1JTaOD<(YZZINbHFN2H#d#4XUCF\LJg\f2RVLLCCN)LDf>C.=P7<W]]7?d3>PZ
K.B1=8\AMWWb\e#BJ2@^\a7c2:IE9\N(Y>8MVc-&_Ae><<9=GHIQMS:DG6#@W,Y0
_)LN-P.Q8,K7f(0)5R-gN0e-YDDYH\L^@=BT_G[/:@+Fe+50Y[N@f,Y4O&RTQ4SG
X/5.d.0:F@O-gR]D&LFe9B)7bHG<LXP?EQ>>BP6S#fXU:G.UO2+(_b@;QYY.TXWI
5cS90b4(@[]=+WY0XW;Tbeb?Peb(S^7K:MBAO0&LIOJed@Yf(67E.B<=V2?BMTZ1
?ZR[J;Bfb>aK,5&E[H/V#c,0Y;FO1APTQ?5d-,[I?PPGN7X9ZgPEH;XP/aQ/7;E+
dbL1FSEge14K3\MQ(A5MA12:GeD4UH)dZIM4M8)fA6COcFC9&L78P?YU)6W&20:@
?,>5XG7J?gFM(#B^Z(Q/-Hag^3IBFQ@&f-.T)FG+#edB_;2]]N_=ZS7-#4MB#e>d
8HNf<U\IOc2Baf;]:(<282AeZR-f;fBgLbE;DUCSX3IKgZCK4V0S(8=2V(6)-+65
=\-76#)?[eX8W?;@7J&8HV[&T:4G\JeK2GBZFcIfS:K@/\WHVN3;S55SdBFe;e#;
J_V7?BdK@TMH&K>Y_a0LLc3OHQE6KWAZ+e8>e_A?LaST1U\aC3-fNR9OdH\ZgWeG
W.D4,<@6SHXV>:<d#Fe+G,fDRH].1GLN/8=3aBaZ/I^JSKN6OZ42#MP[C@](L_Yg
@&AGM_LgN[@GEI329=IQ6d<WHL+9#L18C^bdT-aDf>(5LaNR,YZ3QECg^GT-c[I>
2M09#f/:^2)NA9,\CHSTg=1df&X-ZVgge[@Tg#<HON#JG-?8SVfW+J>BQS+#PD@6
\ENW.-8B,b^Wg?GIW6ePWK#K=O2g:?F&+7(.LTZ,)d>S9,/H=/.8A\TR7(g?SU1L
Y8?K1<74)=b8.J/,6.d13C1/ZWOT+439&AN^/-N\e>;MEQS(\Y4/7\XbIRKLW75F
,^H2aC&f+4&)4U(0c>4dR01W.PPYV]\C(IU8G[3HH;I+cWGDJ\7QV<NVc_DA<:.H
9?4R#_>_W4]?F/dL7S5AN?DXKO/UN>^W.]Q@+OWD276TcDFg><##D6c),W8)Gg_<
]G:/H7V<D]R^>8LgJ]<(e3IF<V8+>2NL?+?<A-I+H=C:^G5W1-0W^f;Kc)a+]/PH
@<W<.[fX4b_O^O9IOJHPX)RNb]<I3KJ4NWAC=^eLVOKP\3(K)]I@>F^FXYN>H]/H
.,d/[66;K0f6T)[:7c_1]We3#2=\WVETSYL<]_S+/Rg(@OD=B(820AS[+X9<J)(@
.(@10T/g=HH[3,b.Y@0HCF<)&J2Y5;B7DNQ.Q&UXFCb2dLK?_F,:))c@5-cIF=e.
dH[A)d,<8X4Z13_3WN>@:19)T12>8bHg?KJ\UWgR[(X#L&X^L4b:2W6SYK8)K&V2
-)V..Eb[;Q4.g6//WPA^CPC#T?Q5MOP,Z4XHHC1+=&W;D4J_<^e>[5e2g_H(f3H[
/Q1[MB,X[<AFA&b20:NRXAO>U4PA9M9\;(>:0bUS4#-dGeN32<V.C_aRMY5QTU#?
D_;?K\6<_RVN=\/]ON;g=J:gKTU]BM^fXaV3-Gb,W6&(\<bZ29?/9K\C:<;gd]Lb
\M2^DAQ+PPM>C_C.0&O36ZGAL)Y@B_>]f/[d=?<?]Ef3VYT4?J_]@W;f<QIH[d3S
56,Pa&)O.-66\6J;e?a#a2)>8G])9JL,bG4I;<ZTA6D5N/e9PYaN-dG[Y?&OU]Y0
XOA?&8-L&F\):U=(63QUbPME&.H?dNf<VKQMW4L#Y9HD7P:DHdW4@D_Q&5G,_5/e
CgP9[?=R4=DAc)YNL,UdGA8-8;AC>1IEcB<2C@?Z;Qg<ST^0]/WUWfg84bgYO/6Z
_NVP/V.RZbL_0@A.3H;Og7J_>Y(9AcX=@H\4#[PZ92LRW&T>A;TI-&ga&b=bU,Ee
3[U#B)=<@98RSeP2#LM7;DXWWWBgHcD:LW#c>IOXC^O[4O]<bMf]B^]gWFH)N2^;
_=39K-Z/YVJ<OL2F8ZGQ4520ca=X&([ZQ9e,UaU=\Wa7)&XOFPJ<9@Y:<<CMPD_<
@I/\\DKV1?HO67ZHGDUGL(00,>5S0FV-Q]c^U9GZ[)8E(1<P?Kg3DZ>@SK?M)OP.
Y+E6Y51N/YAbM.I0FNW30VdNPB/P_WCQFWRR0Tg/YN&)1+IQQ010Y?AcO)W6M^S8
b]KKFPfbeHWS-44ANJ@-0U6H]]M1[BV-Z<gb8;MB3]ZI#RWWNdf@X#9#[GfO]@eE
,#SN7)/2a]2RU&?WPJbB@cHY]PHTY=P[X9a[W==-6=Y)1Z-b8[,M.)UCXGKbgdQV
05X<W=A:4a=_5R>U\JY;UP)6Qa7.P<MEI?S&KT>#a))Og^+P8S[#>S[BV4H=]5/D
(XG/OMAL-G5F-EXU1Ab>EET29-NER:?B3c9UE]#)URfg]VUX6#4gfNUY1cSOR_H,
D=9BgBQHZH\?BbE/]@=U_/;T9:7.KPg&(1<?U:HHQ\4g5>7P+YgKbb?NN<W3+_Z[
.]3IdP(WS[[4\R,Q8Q</Z;ZT=&?O^1HA0KgJ-DFgbQg1S\,N_\SIX&O16@IcHga&
8R)Yf\S3^P1P&g)0=/+FW/^_F([\D7B<R3^_gU:N,3-VTDe.D\Z]a2MKI8,39L>Q
Z[C=H\<D.8<c_26R6a[2g6@,PZ\:P>O_L>-]bHEAbOL/^S=3_VVW/ac0(D9\cW:?
8)/e\ACI_,bABGO>^C?7ffTGCADZ-Pg(Ic/POL7Kg)8\U)2PY9Y0+CN6^U.<<.XG
;9R(N/Y4@[[H0GYG45]]=1(T5f5<MZg6SFFKa\.9=M]^.A7M=06NMZO^^V;3R92Y
7>R^,<L8&G(>>:#9M/gN2\aB[dTObZK;(d/KZNFZCOC^f+2.a2UHR&aBRV)f]=1\
GDKM:/B6<Ja?>C<F^Y;[,:f7\:R^?Y?aTV+@7K/bMdc(1S(F\?Gf==;B[K\79Y9X
0U9GEHBaMb;Zc6dM6VP4XB@ed+_a@HX_&IY(_4=e]MZT1MVKg]>:]>e;UBB[&[a[
fR;:WTc/S)LQWY7UT=-4aOHZ_7Dg2>W1J#13T^f9b[e^fZTMAP+#42eZG[D5K_9&
GH4/_ZCPdY@D1A&-HZCB9LV5b;E)L7/6R4W4W0g]XLRV5fTC#][F_.Ua-X]V(A31
QVBU,:bY8c8[P(RGFKEE2N:/3H)(3,4Eg&HgF#0\.03<^;A1T)R&Y28Y#a_3f^ZL
.RaE>[:BXJPE[UeN.<#NN>OJAV5_6&fdPdF@HJ\DO/VRN=2#.RdE97>K[K;+O<O>
=TBHAZVP6SJVFS-:F<-[#YeZCKF]0Vb#K>Z)O[bCG8bV8b/4#FfY_O;_UYXgU)bX
bD=(G#,&98\[BBR8dU1c>/#_]WO+CVbH;MV36FQJ(MC+aID=E(ZEJ^AL@S-HH=)(
fQ#_9ae4Q&fIbN?:BcONV^]gUWR:/0?/>C5=)SZRHY7VAU;f7G[PELM<\]PQ2Y6T
WVY/)[H+G?+YVY_=5S4ZHZ+US0UgM\7=22NJUg7VJ?L./L<OccOQMGUSg/MW&0^K
]F916]D6F20cM-YS@OTfX0,OZPZY(P]>?PDMK/X:P]T0,ATG>MK\M2gWL=E^W,CQ
DRX@Tc50I^>G]^6NKfUTA]7T7_8U[[RD4IfWa+J1e,GcOKc/MTQN>9a.@L,F7-I>
DLI36b-.K;bKVMU@XJY+\0cZ[geD,/.)][/K1,&YHaDDRDI)eK3CVb0He]CF_J(#
NPZI)ddd@O7,CAe+/+6;+)FaP>]YY0A-?.OJ1VdV_T#O20dWP00DZg6)OY<M5K1_
-3.1J75@8G5bA,NDJP-[]RE1.f?9^4SFEIH7RN+^/L[+^.IaZcce1);_cDLK&M)S
a9Z;21VNAAIN9bV.7We3P2c(eN(5E=BM/6&SgecEDFCdI4C\FW@Zd\6TLQ6&<J(6
FfSYg/f69^4Ed5W8MFE[MMS[=B4/-G,eT5\;?4?;?L(;B,280A,0(?CE;R\f3?[2
3_DHDcad1205dDH9\5<&d;J60]0_&F^5GPT9E=aScB;&1g2V>=dY>b9V/_Lf0Af\
O_/A]HaLIa15:YP-8ZG6fW3<<^5D_3Z-F>ECLOK_>P:,;9VQPJ&D<X9Ka;I+ZW)g
U_9<.=/EG>7R)Q5&F)30b8Z).3R@T1bFUYNAM1.U1NUebTc>?^(+P47.ZaI8b/c>
,M;.^(+EO,ZaP6e,Xb)6b[>7#g7>P8HG2O?\,(H1BC0Q?;89A6+,17Z(&LG6gE6G
2&5bQE:6E?GC1^;>VV16VH6NDV=cS?DZP)C4PbOgJ\PCdJf1FD4E8:7Y[aDG8aL#
W&eC=K(W1FPf9c>TYIUM3-U=;]MV/ADRB^R<-V?-g+_YZ.-FTV386EIddW1GRDPg
8g+McJ0RB?/;\@;6\Ue^;SAaBNHWM[,42ZBQ#77V3?8L?W->=[CF=<^U8gf:gSZ,
)B<^^#WJ5NZWd@^aPQeTI@VaA(PFQeB&Fe1^L)>QYY88J6DeeM_dJN,?.G-IITVI
IHV)ffS>Q09]#K0DMV5,a<JOAZ2QZ@FV#L][d>-][4>K/c8f4GA^-0N&70B#-TW:
..GLF^:^XRH3@Q2TR(cI1c,08S02.PU;<(&_fcD?]/1F9eG[c<[6F1H^=@(XF7)[
O?#LWTY1PP;\V+<+,;a5@f5GL)DD/LMS(.\LcFY[Qg^XQ>/b_e/LB[=F>HX^ee\b
TY^][W2P<Z)DbP]E35DSb0;TMf5..46N?DU2SK?TT:0Hf^1/GG0O4J5_6;f^\:6J
])9.2Z;/>0++-URR5KKW]bUU+UC[_8ZM&#ASN\.=8<Nd@#1eL=eLGV7_1YIXfF^N
LOL7#G(e:cW)Q1F,_HYXN:bG4A@WFH.gNILX]-f.)5+WAJT&a;/IR8/:/68>5#CT
IV<F[P?DHf.cV77?0LC,IA/>:E3aNW)R7<7#CSfM0G?]QB38LJDL^;L&5gd&X?aG
31W=5?Eg.07-KTO.H)PVFV41N0UMebI#cffK(WdQ_ZdR9e2eI4+8bc]d/_ARR>ZU
]6CX?PBI1P:>&V-=RC:ETH16]\<BD=/bGCc^CL?ZVZF;<W;7<CGK/^;FMa.UVEP&
_]EV\.[Ve)S]gfYZbC]@23RAH-[V@[aT_bZ9)[W.d;:6GXg0+ZL2c^QY&2gAEZ(U
R[-X@dUFbC;c+0XT5FRB+WT(d0_g3Jb_7\#cH^NM<T=-#:TC9@#NSAA^>EPM-AC_
?BN=3a&?ZKVIbfQaeNOE<_[9U]55<P>C<::<3Q?]SQ._SSY=>;P54I^?\e_QDXLB
46T4dF62b.&[g@CX#B?aNNE7=/[?8=_\)>_WESNdJT]O?>AV9XED?.Wd8.Y:dG(R
U):QO]:N4TKW+Yb:O=Y>L7FTJESZde+97-aJF;eMdWOBc)JC55?;(8:3(f1[JP/M
_AWJd13@6MWB/.4GY^bSJ@>_b9BYM/7BOA/5#()&:5D9F+>P2=IgNKd)L-.4XNdA
_ZYDd9^2=F[@S4@1F&_X+B2S9P&V,R@8S1&NTV^O8O]X(5[H\;9<&/^N?MTXg@HZ
]8Y45(N+CV-LV]G=F<^E<TG+#QPX0M60bg-A5geRIJZb\^C],\Je+2]D28I#>^1M
\b66ZAD_O-,]RUXT?6YIH<UJb8=U1;)#FY3HH5>10g]e]5B2:_\3K<Y&0U\],6L<
4ZQ?ODMa()1N,I<FCOD;IR6>gIL[ZTS:0V)c[+5[PN)S>E\UP3NQdeM,)FSZ3(Cg
SB2X^KR&0cYOXG>ZSd;T\^9[_VaY@IDAUK=&JC/FXYU<4U1J8e5DD<6SO=&0YM&<
Z[.H;eVe]g&/M3B189L96b,\bGQ]OXD6XL7WLOMdCBU?Y)KLXceJS(6D[7V>^=Nf
>b-;@]fX&F7g5SKWG>>#EA,QTN2YBT&UU^PK4UCJbd(+OUN1;[YI@O@,U@63\,#K
>eHbI0O(NbX+V+FbUc[;+3OCO8;=IbAL5ZTM.WQNKB-O\RE\U8gUF\D^4&WE3R;R
Z_A-TC/@U),KZ)eYW5Y08>8I&).ZF#D^N)MXLN;6K/aXS2)cL5G>J_0C;RMFW#P)
\_;TUX>O5?>1QaTY1F4&=PGV>Y85)D8RYX&c9Q2S]IO-O&VH547DY<f=@ZI>Y&cB
g0]a7GdM>3T(97YK#A)_DJ_<)XP-cdDTHG<]>DT;X,#+W@f7b(37#gbGW_7[4S4;
]5]=VEI9&REX]5:;>>ZF2@;40HP0W^.H@5DT,/.DL6,J^EV&.MYdE;]Q2<(g=DOA
6UW-E9fPC0^2gAHF.Z2P;?MF>AR//^7C.N=^22<0?CIQQE]4,<DAL@1_3,(Ja9PL
gC&8AX5::J9fAbY:dB@[U/IW?A>8NZ-@:JFN,d(4^[Z-UN8_1aZ6Bf,MA/VEX7OK
;Q:R7S(&)FEa<M[=2gK_-^GF[@M6g91898QZ\[/C78bU>6eGd7EeacdC:]bWA#M&
Q8BRJcNPN@,42Og#/c2e#,O1:e7TVO>XJ[H<DFLJWf>7N:MDBCR->,^0S4#@?.ef
@,;ET=DWJF&5L3(U(;#T\B(G2>4X;;L5LKS=edOUKF&;EAb-?AaAG3_f=S/=YUQH
HY>J&Ec;5F)<-.;aPcHJ)=[++^A,T@Ad#DA5bZTC<[agQ+aG#]V72Q2SS0\_5Pc=
PJ[L_Q^&HB=FC5N-2VD=Y5cc1)&7F7M8W[&K.37H5]f4NZ&?0339G4O]B7NS&##Y
a.UHO-I?910VFQ^]a(.KMO2HN3JJ2&FQ(]+c&-Q1YQ>_d+\6?[^8a&H3^O-R-0G+
+g<Y[.(CO?9M;EC[:@2ZPK142\5NR2_(d=gDZ[G=JaTWe/A9J)ZDa+7=Cgd2ESS:
MP]AUac3aF<V.EeOU[YaNU]GTM[;X&:8&Ag)=QA#@06+IgEI&fUMIbETDCZADbD&
:CK;><DdK?H4d?8Y+5T?R;?J_DBd]JYLbK3.)Q.\)WB&#McZ-00bfIV?DS05[#?(
ZOaVY;7^A:L:OcU6M32^6,&SKF_DRP1&D51F+67:HNGJX)4H[Q<14P:_/c(,Nc]Z
F\<c2Fg//6#:?3e;5SEU<<L\AAbCOVE9\aNV6?B26[ZHRR15&<6K?W#=77_?M.KD
_LQ0F4LIGX-aUgMPg8[a)]<3:DPADD-=AAY-7D5[M@L;X.+.Z7bQLP/;gc:N28M.
a8Hfb-?@d[f.Z87JZg?HJZNE_LWHcA<2TRNRKSRG<FdW/IKYXX.D:DTc5::L0Z\J
+NfEF8,T)0[SN>+>3]T8K+,@BS<E:-K1?>,JD[1-aQ2:=fF]&cX=d04J=@HU+H.^
RO8;2\bEB<+4<aD>=SKEC;JW].fe=LWG(;YAT)_4;GG1/U+&@=7,+G(9(TgKc90K
;=Y1@D@..V71Zg<N@fQJ69@/gdR>g0Ob26)KX5>-,)-=QG[]9_J,Wa2K&.5Bg7S4
;LB;9;SUP_6D+V.fV=_NJ4eL\_B)N<W?(g;HS,K@>-_=)A)PbY+9bK4dVF&->G=.
OC[<a6dKg#87b=B#DJc6a?1.ASIP;&#^K,CV<fC;2MbK[aBIe2:b5#].C/O\:7K5
#_/d6V)EcP]aL0XZYXQ8CP<a>AGB.5S.,9eO65:]KaCR?^]CgJQ>[YeB,WZeOC/g
)RMd>RIgJIKd[F#;(G_R=E.K04-#0R,[0MJga?><8@9gJ03-\1#EPPbVHg)M/g/E
]MA+2V0P<F6UX7DSd3A8Q-M:7W,\gJA(:L@26_>b-KZ:IZSfSXf#:HPC,ML6,dI-
Q?d=OO)3(f&b:aO7Z((36/M55f@/M@27>@=JSRO?;Q5S2J:OZM)3Df]>C+;RC^Q?
+-3,?,P^U2[;7&-NM;J(9-]6D18#BD19ECF72(\gHM,aV_JZIQ:Y\I?N(C<YL.]O
IFFPZGF#dRDaUT+<)=S;Be[HA)+f053SI\[CdI4Z],CJA2[@\Vb.>,c4Yb2JIO/O
F8_H7-<d,d_.TLa5T0cEHbQ3-.a]F99(XgDD;D:)X,:ac1UC=-@Va@P79=,\\4P.
L1C-IfSQ,/?BU&2@cS6K+T1=BHe5b\,LO)P;6>&/:..I4gT4\0>LM9G=2R6HA.c0
a(>:)#RUI\IPVH)05;Ec0/1G-gY:X^F0BCc.P2OO^9/.MJV3Nf:+E&@Mdf_VL@(J
6YQPDO_586G#5F?d@DK)4^V,_aNW^2Z/<-0g@3R_8D&):.K?PQ:2a/LdHb66,VI_
b8<A=>\B>I[8DJ1]NE55,fUNQY.a>EP&#<W?,-)HN&ILR22bE,OcT+,BUQ+3.CCZ
5K,SC.LM=,9\O8CCO,E3FSN/UO>6Ja\TOPA.f7>6J@T5eDeG\XBHJAZIIdFR[SIS
4DL&-/391AX\IBLXfC<E=[PL8N/eegZf>Z>R:NRFVUWL^S\,-SG>CLQ2cH/OI:&.
/U\1;#4\e,@1f#b;&YWMDfRK89O.CGMIITN(e39I&C(cQfR>Vb=E1/:G.+<\Tb?C
g..#8MH0)T^=VOS^gQL^4NRPZdFN)8QHBa]ZO733;3&H3af3J?IK6&?NUg)=8R:N
^D7:(9:GNf+F#ZU:+9TBaR[/A\0(V/@\(YFYb5I?d:#:<dM^YWa@.-&5.1HeJO2Q
da\f]?QVHJ-TZfX1Jd]@#gM<6W7GS.+-K)1d62aV,.#JT8096ZREHVVSAaSbEKN8
L\+Na3HGae7L_,G435fB(/If@7HF2M0,d[A0YLM9^0<fJI^]1R4?TSU:2c@42bAW
Z/PKf.9AS=C5KaLXWJ_@F;d\_8Fa,<K)KK6MEIPS026,4^fL)\VTBR0IM.-<Z+:^
M5.g3M]7#YJ.H-H^B^C3aZbIW:g\]>7[2I>,Qf3=>6:=eYD.6:<5@fK5b_]K_abY
EP4W:f[g&MMFd7\EV/d1EGL[><c;Xb9C[1=32MBH2:R,7aQ=>Jc?O7K4^FZW?\>K
6SI;_YDO>Q5?.:91E=?a&F)^^Y6De4a-KZ&,gZGc>\O.Ec&EB<U[aI[QX]JcD\A0
DG8@GO3\2WA]WI09e:WJ[W,^?,/X2(/4RbAB9\bfM-[T7g@ND9e7FSJgUX;(T_MR
X)@UEf8_SCJI;[DEL=L@F&)=2gBbKG+-IJB#gaCB1SH8C+;>\/FfH[YLB,<P0RY8
,I1/=Ed\@IC4#fWBYN;Z3Q7)DWc#23W,[f;O;T6FG.ZfQW4\62XKV+\5(\@7WG^V
;_^C/Zg04^[E:.<@a=?T)cQSM:=TVXJfRG(\QdNT5b9-WPRMg\I9c;b^b#/O:+=H
GYJD&^YRFI5577(?(?1VcD0<S(TGS;R#V&[e?][VIfB-fJ0UD/\WK)K??GTI.==U
WFP[J@g/JO[2#N:Q6J)Y92+a@XGGI.cC-eN9X.QC_7WaG:_.[T2ZE[:gcA\BVN0,
=2H<^?VC;.^gVPIg)@1TXC\OVX(O5FbWL8BFf2V>,260H)5GbegE[=<dTBL,&b5(
\JX;OFQ:Ga)XD:/Q<;.NV4E<U:]3>;?9;XY)dKNPAT_GP.ZPNF-T>=(3T>=C)a3M
KPFL82S9MI+DC=X\.DcCZYQ>OFXCc333MV8C:9dW_ZOYJC,Ua2DO+_(,)<923J:f
=B]AYOgN]3B;[[NcVUB+/bZ=C.#M060WEEEU]Kd\aV,[9>/EGY4aDXIHRGU;cFW=
^9]OTJ()Df&fTCgOJ7]O2c,RJIBDVF\KMC_#>9D]I._EQ,M.]W8+@=P_Sd94e<G0
AHA<?Fgc6+[-^.[6(FY#[/?3F#M&YE89@TAYV_f>4L=[55LL)3ZdIaa,X#I7YQ&E
3[A-cJQ^1QgWW[X_<JQ?1F.1^=6GVG/U2e88^M#5QRZ_W@b(-XbJYb:)?[cN28L1
F[W&BV[a_V,V08_G^\&ba/gR89&9<O/W?@4NV:+GT7A2SKOY3?f&7]B4WED+@5GT
Q^a8#YIa508&Y[FJBaW(aH.369_5<;+Z,EU9BcM4eaCP-9)P9.d/fX)XbD627U#N
#-__?,0Wc:J7BBR[WDfR5aKDLH4,c@DFOTXS5L-/N27UEQY\fE3Q:<9>&FfKAA)O
(49^Hd/ZeQ3+BX4GP#E^OR3<>eSM17;aD_aE+.&<].[6L6M31c#M5F)P2^Y/ba71
:?R61D94J2=_>.X4Za.Uf:>7@&R[DJ:]0_JS:DE\a\[M)TL/^WD1DZQTM9K7dM/\
,CS7ZLTHD64cbadfcST7@52R)NZU#FWHL;R3EH4=fH9YEeDCUb@9?/#Z5(1OD0KX
[H/d-53Ga&SL>E7&WPX^5R278\9<B)AeXMd;NE??OdH&X<FKWOH;A^+Y)UR:?e0O
1X_0Eg?19\;6J[b5cK<)EQ]Mb?:_S[b96W<A#;DaK7dXA?6JE;Wd_[8:c58@dNac
.0FV3<:]AN.W]JN4>aJT,O#S)O[fD_,E5>IBLbRPQ-S-F1YR.aVX=a]R3899>NZd
f@QX/8G1e6TDX5)Z0Q6J\5^UN+K+C;@.4Labd^M\feR8B@#/^e,TN]fa>0QG^Q)>
_8TXKc0ba&<UbPI4,R;::KN//FA-a/LB,L&R1[&K&63OML6H(5AAIg_,7GFXTT>:
/bZA]aU^<T<1U/GP250O;U[I2GOIS:4M75X3@8>e>gV8W7DM-P+G&TKC@A/FA_\9
7K)Z4E\e[+@H5a1c\eZD-GK+98<(V.)3B7X&CG@A=_0[</#Z[BQ3c>UV84@bV.g[
EY9#]Re]0^.(^T:P-A.GM)aLC2b_5X;RJJegc<\_R9R@:P\WfDKd2Va,a5@_ENT;
S1a#3Q](I5>IDM/8ROXWc.Ja9e;0@NZ<ad6--<[RDLNIKX5H^:S,)]aS@^^R2_)(
LENTW][FLgS?d&DE+/#ERYVR9G]J1W+,I6D+30.OH<-T_IF&3_cL:/LA?M0S85[C
S(PNL>FU/@C#.b9+e_a;e3HS_E[/.TK7SX>/DI,:J):-,7K\gdQPF],+?\Ba8=I9
3d0a^OAcOM3M\QGb=U8Q.LeS/YDd6bQ.<K9VAg_Yf,RLJ8ZKZXF5;c?,=)WWC5@)
@/6R@YE2SUV6(gLU(Kg+G7TAV&;W&>]1I5NN5DFOEQO>bOa(6@#f=Ae);J,TJA@S
:WN,Gc#a32_g6#0OMSW)2K5D+S1PJF[;=U(UD53;?d^0<RF&MS3NX7F_)feg/UZK
I\\91E_b>BXSd\SX0C@b/O^CagQ7:>E(AK:(=4P6YT1&Xc/&67F-WYUc,C3GX7,-
0;F#))[aJ+-T+7W/]99][9X@0LN-_4D6T;\A[fU4X.5@^#YX6fLD5CF;,dVLe7]]
dSe^25I/AX^E&8=19Le0F/OQ^F9b#J;NgMDNBA6Wc6LOb?,S4F:EPO872d2L_M3V
>/1;K6]cE<&I;FI5NBIg66eUV+AZ\(d=\+cZV>6PW6FKVEaSW@R@/D9bKb=3K0eV
B?#;IfG[3aC0?bD:\[0TL3afW]Q=4@b@6GH>TIX&Q45b9#C2683,W#UBN@3H7[][
2-+7QVX#+BW(0eOS6<BLM31+;g,SV7g\Y<AM+>8P0eW7a(4I)@Yc#F=MK3B+Q=68
([>>0Q8Q\\N4B99NZC.)-DGVf/@QWZMK/I8DSLEI@;P<fX^2@S#6TKR7LV_Ka^?A
F&&GX28EV=UPQ1+7[BCb?2[_11OEae<7?;)_P9OfK&QV4G7M?7/;XJO/+;SD2=bR
[].JAJXfR=+:A\@(HF+0@g2LL/K1OE?4XLIQ476OZYG-7_(cE^JLcNS(:3^]OfMX
-J])</^JCG_R-e[eK^C3[.[F3=_PAWNYPZ_>+7HF0Mef7+JIZS@H6/?WJI_0MRFD
C:@O1,7&^.[<Ufe7/^J8F\I88OdG>\],O]28A4e-[3#(QPdQd-#J7>a5&O)T8MeE
7^#f-<OX/1.eUR?M>[=YO-4SL5a,C+V0@^PeE,08e_5+BcH.>?[Y87CS46NCJ^#e
E2E:S-TgZ&S4BcgW:U?IJ,ZN56Vb9d+I=6/6NU,;)g1\MO9\b?;O((/d1)0D)4^:
(45,g6J^#<F>R10J/PG+KJME>GF\Z&Ya7A_4e(NXFQX[<fZaf8#F\P^g73FBJ<A(
G5/+_YcNT>=K]3:DIR68FAS)DVH@+bCZgbdP&]:OY]QG,YZD>SeR-gX<Y^e(:f47
R><GBgHK=XRO^WGTKFSL-<9UW&?N[AI-<FK/#3&+cKR=<d?0?E55SLMG?UAAdPOS
Xa@/F4:F>e/=)X_gZ1a?S).:4W(@?;G4&T+K5(5:\7BM/cV]:Q)c=,9AXK?F?@d@
9feM6f>]PJ[=6JQT8O;<@Yg2Y()7?QM=cWPc+>.T]]W>,U:3S9M?^[ecV-6e8N>E
H(S(J]5Y7-&OY?[\UI/7L/_JAQ7IbC9NNT0UaRb++7_E(QTg[AK&&_NWM(TNWMBN
+KPOYMgF?8DLVMV/^>^804]aG-fgQOSC:b=FNV\)^g9MZ0S5#B/e5R@<&E^=)C&2
=://YK03?YMTTE.Gb-MYb/?.RBcO^NJL43f_M8HF>1#^>.,0JNB=)LS1f[7KZX._
O\:X9.1aQILRA5G1[Yd<YU5ffJg?_AC.(0=Vb@db@d<^T18=HUg8MKSCH^;eW7AO
AdGc&MF+5?I_GM/=,\@0H-gAgI(,3NF<XL=0bgf=PXe]ddLNdTSO::P>=G9(f5(c
b-]H)OP&9N&ZE/]2dUFJUJE8,Q)F<#-NPV>]IH_Rd5)cO?ZQ2f+/KS6[R#6ZSXA[
]SHNH6#eLQR:2]0DHR+W]DDM,73MIJga\T(=GGA6\2QDZ+&@-PI=^H<P;8^F0HG+
a:=J+b(BX4CZ-7/?\=@\JD^IT.(U^LQNWE:JYB525TM2eN<2UCX<+@)W=,(P22Wb
Y@D6?g-QBA>FTK=@T.UN-:-;(6I.IP&>\eSgXNRfQEVJc;)TE)0IPEK?<-IZX>9P
6IR_PZgS,#0\d#CCBUDf<e13X+-<;6=O^&;-@QWIL8:A7PLP-L8D#[Y1M7E3WY13
g(8f4K;C5\O88_T1Yd)SEU>Q,-X[bPXg-_:aR;6E]?QfGF^Z?G0/V].e7PVNHe,U
K;3.G][Dd=UX9.>P(=#]#Ee>@\FaI@g;cA.GcUUYgL@E-c(+E[,0EZ>4.R1=&:HW
NT])2?UUYb&2WgZ1^?2\?,>#=D[TDE9DfbT,1aYRV6J+]68Q_SR+@AMM7QCGP(KX
/+9>FL<OH&5U?SeV0_4b_PQg&EX?c3>P_T[N=C=(JA@#L:,ZY?DaN:a\IWB-K/DK
B+8aFI,4/)A.HX5>TSBa<Ec=?@(\8D8S1@\UY^bWFY4(:B>\Uf;0HSBY&d?UH@TL
)=SK(4Qg>Yd,51dH<=\>,e0,S?OH4&;eaM4PXPIcA>((F+E.7BRd4[]<D<6:&S]8
JQ<aeOaPZ3bT:aZ)Og5+3RV.P1;Y>NJ.S6Z5(Y=IHE>8(8F::9SGYI>Te>c\Z2/7
>IP#9I1eIT?<4.6FaWRH=6.Z<=;Of4W(AIDL)&.Z:GPATQDb5aNSd-@D)(@f#<ET
+b8HP2VDDV3U3<UA>UPB)[[2_BfZf+:0Q@+d:FD43/>PNZR(GH5Kf4;^a5Ba@NK?
#8DWWTU@e4:9DUY1e,PY7;Xd021KY#(?g5CWL<aSZ0<AQ[4JR0F=360]S^N2fJCb
MM0XT\09/aW>+e=]YUP(2a\2LO3SDD#^.2>V&77,J=GKaaK5VPYCD99DgSYR[CUF
c,BFR/^1((6(VC4JDWgZ-9KQ1>,^U=(NNNc_#-K+e4aG5W=JN].HF8&E,=e_#>MI
MM#4fRZa5S#W8TcN-S+YL6Nc_>B<A=d9S@5?#fJP;9-Q&0fbT42X8@J]C8D=FDE@
.5[AT69,#DaF1.^+V.=1XfFTC@.^DY&5A4F:Xb=b6GD&]B],X:^^;NJ>&cS<^a6P
XP)>+d?C1-S@?M5QD.7LV@SI+-29=0f-TR#MFO7)32_<OM^=4\3)(B<4GQ9G[>7Q
aUTbgFMNf8X1DSb(JGNLN2CJ[+a^cYXY)Q)UEO\,cfP+GdXDQE6;J>W5\C8A717J
;&b398c@V4\6NJ#N>4SJLZ^>8TOR#<4QN8D@JW0J8GMV8__RH_f=@#fSgG5[W8V-
\R+5=7AG8Pd>\b_e#DWNU7Md:ZR+/RZ:FJSH^:LF8VI@B70db1XURQaIJL]=Ted[
Wc8PRW<?Ab)6=WQfR])>f8K6LK3[^G<BNeg)#ZYRI=UQ;Z6AE1G]a)8b^G5F_<GU
.>3JZ3-Hd+AT:323<83(N5UCgN_ec\^Wb;YaV[P9OcU.@4EA?C/5C1V^1Wg\.\H@
VU,_ZG>?7RZV^D0CZ?7LE3I;>^3G[H#6INV?)M31#8e[HUD]I=8^_D_B/&A]DAIN
>(@[=VV[(0+fGWXAS[LB@[4Vb@7RX-#Ka/10A+bME=UDSGJ8U9@6G@b2C,IQMKT_
f0,U7ZP^6]O>.487V96f2O?8--K2UR;<EO/=,Q?-)cAe)1K6_6^LB:KR4>Z^?8-5
>R_R^P;>L=J8UgIQH,;4,OM@1G-A]F;J.4b+Tff,@>=:K>dSOUFeKN:7;D@/AVa&
)?QQ\G\c(P;3=HERGBNE]L@Vbg4/Q<f1>9(bU\e9#OgHITBY5gK=KS:A\X\@W?+#
f^#8TFGfD.gWJ/6a0bQ=I;O@[R>EK8_ce73J\dG(UPDMT15+?cJ<f2=AU\5/#<#e
Kf/-3dR.43#M(V[I5VV5_aWN[OXVZ4@L;+&9D?>D2MG(0B=K2HD49]HIJ+D0cL@G
Mc:J]W@Z9^5,?b55M(DESQ,0-DKXSY0XWQT528==A,<a#>bb-=KA-^.UaGYe-3ag
>6KH8dIcX]dXY7-b\[.S3]Ga8PV5M,b,?GS(KA@47EZ>^/[1KCW#T,VKDZ4fVb?^
O1W.f?IW/0Yg#H#(^=VJ8[R3f?YK6+C>+2(ac_[812RF>UbPbZNQJ?S_6N+DH/90
M&1X7IQPPH3^64SdCVW@<B<H1X_4,,V/H4S2>:_NF-F+<c\VX+C;0=E3\?7LH9c:
YQ#Ned?^bYZZ1<bcM\XC:/;.0bdJa0]W]-Ned8G\)>NVRONRg,\YTK.7I&1&;8T-
1M@<0@_K#9#\T9N=NbTaK8#00[.AAKUYU3Mf5Xg[:^26(BYL1+b@8cf_/ZLSLKBL
]V7;-@]Q&3bBJ^IBZJGOaJK9C,2=0FO>g#AJGCUTAMKX).5EAa/gVSY:J5=U:X5A
3LV[^9[bD)Z2.c#AS[<We6)R&0-Yb(_H9&KR]dB<MNSC&MZ^G8S@SWf4==E41aD/
aN<0S/2O>(O@,D9B^O&?6K&)ELWJQL(ge/^1)?WI]KY.RbC5BJ/NB]GU2;NVU0W2
JZ-Y9[Z,B?f7))#C;gP@7eH8M[)7RZ:B<&d]ZVEYGII2[9=gM^,KV/8X[?:)NRG#
5d,JUC?^Z(YF+6K)EY33WFN(FU&CW;VE0AgXKFaN@Z;)5F]EM\IJQ@G+e>,V<GAd
DENV74QY-:AW2V]ZY,G+O&\LG#H(IbR-[@<gH8)VdaRLc^(1:EA=R1_T6#^7fKM\
eNAOF8>S-KKag:Z0=c<:T9K0dC:LGIH>1;LKaY)E7bKD>>8/c25]1dL#:_=+<6,f
1&4aLB/1=,ZM+fO=dec+IX_1_1R18Lc(EYQR_CURL.^EfQ8;#LT=A21&#7-e?([+
UZ2><(2TYQ(?JMJ55b,EH;EN-[)?D3+LT4Keef\Na?a^Q?)YQfAPRMJ17gLI#N=e
aA?.aKDDZAKE\\/9HD0#MLG]X/3J9YaADCK5IURDZ[A-^HFH](08C+B49.FHeM]W
=P8#.7V_HGNf^3C86fcUfG22E_KgJ[E[?b2@+8Q;U]E5e4(8[?9NPEXUA+(?&;Ad
;b5N67/B57Q4AOV)C+::7I1V-?)8:C^5gcG:71-@7EXc56H#9O_X/DAC\C4e16-Y
1HH_-V<Z?b^]XT_5bXTcUe:2A,[O<W[E.<0@8)CS50QM58g0aVW&Qd7&T_E7,6Jb
U=A_QN=QcGcTfWI5f=\[I]R-=BdPcK=-GG\MI>UbPR<a>PDXGR50\Q/3>#@&N6B(
=_NL0./Gd#(]C5ZVMX#CW()EU5P<T[4F+=]Y^WLe_[aI<SH8OF2dO5[010g7e+\K
[9--\3FZ6<1DIL#\+#f&?J;&W01cI4,bIA2<,<c:&,_<DFQe.:5@Ce^a4;E2HV<g
&/g2ESP,dX=AQW(e8cO4LWY;0MHSd:Pe:0cGg7SG3?C-.#_?d/35D)0Q+\(;07fP
Q5,d=/V?,FM>WZOMEPER]IBI5RL0G-@S6JcXPQ++5Oe54_#McY4;/B7eI&CWG?U4
@K=A)9>,_&@X#@LKCT3TS[f>L6V,-H]gFBNWSYV.2egT+J[GG(A973TZ/eZeXG9g
I^d.\NGE2UT3;?]DL73a&@1=bIJB+6DFF&5f^542eO)(Kdg[@2bR(T3U3MCd0TdA
.&9Z+;+.0bggZ)O3Ue/@&ZA(AGY2^[35>aX:DX(+g;)6:aSR)_LODJTTeV856d(-
BdU\P]3LacC#Fg.>aWJ+DY?)1NUVPQGc@EaEI_-/<:LLK_&_R<C,L2/+0]gSf0X/
a0UZR2=eRGDYR<U,4fCf=S&\&+:.c6U+QQS8O@CW+PQF\MY=(fBG<a9I52N2LI^B
OH(.W[eBbDRR7R9\9:30,5WBRcO#B0152QY[^]GMZVL6UgB+I.>M>B4c.eFIaA]W
/(LYU&D29D5<A\b@?,VHQPR;A.HQR::C@KML5/]Q8R71c-&0U]-O#PC/^3#93TS-
5P8\Q\N&5JYW0D3H^,8Tg3c1aK(_TZGddHMRO&g=DP2WaIfWDUI\CceJ;NCPNJaR
NfO:g+N?.GC.Na?BZ-D\]e^99]?F2dMCWRKfQHg,\@-E,MP.e06??U#KBg(gR7RN
Q9PB-LcU[BE@L>G2H:7OJ+(f)/95/dFJK:RQP^:JEA>efJSMP/A/SD6/Z7W]Z;(9
/IV)fU.75>30]_>MeTg205(-IV&^BB[-P=^]<9=cK&6T(g#I<YLa?;,JB9b,\V^6
;>H8C@1Ac<dIQb3G0,-SPT1fF6ae:;JI>^=ac/JeXA^9<JW,=]\Y\CN?(M0BFM5a
NBNA/>IbU-I30R]-VVH/1=9\e792&Q<4YVJE_VPU7gOG^Z@9P>X9NTKFU/Ng\,H4
Mc=FA>&CE1=9Ee@?C(/ZH12BY7@MW(WWZa/2L-6=RD9AZ.d+?A]SaZ]D0B6RLJ4&
4VRB?F[2,-R&6=STV[a50L_<J-,K.4K,=.[H7:b>Fg/YTKGK5?U201TK\F@)FLLb
45F2L&I70Z4f<2dD27DXM(3G<7AK/R^R>-UdL=gaS3:#,Q@K=Ob0NfL;Z]SfA-=a
74/,>3_9RbXYLZ?W\?VGg=M?&g6K+98>\^gN=3,@N&VS\S^.Q=R\6^HK8C329a4M
e@Y<aK(3@+2;#<[IM>&,/7Y=(SC5cKa[U(U#VO8ZK1JL87-,F[:2a1<eA,^@gSVa
K.ccO4^Od7S&9e&M,+7MQb1<[(C<[^>R4SC^.+N\4TR07GZ4HK7LV-aHb>>O0Q@W
+TXA,gaRN?.0XM8N6c[X&]C#SIJ?MK8-aW/,[dfZGLR)@>^+RW\2+F>AEG\0SRaN
>6?1X/=TCC#_B\,9#VWcbg\G;=Maf^4aA3/8gW>RgW?0\3+Q4.OG3KddI32<b9W-
<SX&>ceJ.<ObEKAVO7>)^+Nc]4K3d+ZAT4X0EA7dZ3#CKL?,YM=1_b.]D3[#MW0Y
c4Q5d0SSPNbKQQLJg]W&6UH@?8<TUSd@]DSd\MWC(&BM5208HEc7)0BGM5ISDKa1
gSbI3=GcF4P._)a\eV(RT5#W)CWQBf:R/.RH<DGH4WZRKF1-YTd;Z8CHc78/DOC2
OG3E2](ZCW=3T[S^KF2>7MSS^\?PLG=L9(3A>L_G+F3a?>E&<V5Zc/7fC4H:NI[7
bYAXMf_T:^856F;O1+Uf1>+FH@BM2E/HS61YNXeKY/),-7RUJOA1@OLCDF+ARUJ_
@J?CZC5VeJ701b/H/VBYZ0)AAB6N5)QI6BK\/_6A6D1#4YV/@D+<X(+R5^K=6Ca=
a79&4g0S=FY#AgLaIB:S<J[)<=EISP\8[O2;QFS+dUHXcG0dCXC2JD1G:<e#4#=3
QB6W-Pc^P=eIe<cFU[BCdS#c>T3/=M[dYDI8U=[c=3PD3];MSJ\RHIPA:;KXHRU#
R0M:eP)(eXQ8\cQE#]F6VK=XHX?^,CZ82,NT)PG13Sg=>P\YX8Z++=X:A6<b0ALF
2F/&dJ3Q/gP_3\ED:H1f8N=&GU0BGHZeMe(_b]SHDQES]b:aNY=V0Qc_6OC5=QN<
MeJb0+5+]4V1+@615Z)8UaU1\;g\\M\Y1I:RS+.]B?R,bNL[e+&DC)5eT?9)b8.K
UWTW(@6,IXW1YNIW[Va<Z<17bVR,_D,]=5Me,P2_bXOE-&Z.^5)@dETc,,5ef@Pd
?F9WB6Fe&)41La<7.@FB),&-4/#Q]49QfO>.OLLgP;MMS#F;#:?045^#ZT\.W;U6
;97/)WbQQ/R.<N()C-PKd1YZ>X[E#TDWROD<^A>bF#F(#9e?a@fU_cFDYa?..T)7
Q((DcTDJ@INHS&KIN76&AY@./]]L]SKQd@=VaJI<H)c5gBg+SN;<<492W.cRZ#HO
J@4LWI#We^G9PTOATAaUGEN@/A.aaFKF.T-[O>=Y6FZSO(9PFdWfP5]_9I^g)2ZQ
\_CBBf=+,L[HJg+XXf=e11Nc51]DGM)=ZV6VT]d/68/We8BaEP.DIZOAIA,S#W81
UdME@GDLUWDLH1C1HdV)D,WaLeOD&<L_f-ZKbOH+;e]&K/<\#=H8+63+LM,U@5G6
C+/8#.>FF)E,<2Q;K(#>0B+;PE(9<?>P4eW4CZEIJKNN.K\:,O2UWNWeT?9[<=D2
Y@YCc8)b4A-<ZP-C&I)_D]4I^<Z07/ObN/#[,[Q7)#JXG7S&:=<KQ71>C&W/1RIM
CP&&Pg;4^H2Ve]([W6g)P1-f<\_3Gdg8/P@GZW]F]E/\6^RNJ<+EOHdYHbU/WPd_
+;T6f+UARZ(I07/P+HcSC_1<.?+C.)N&:Q2SR,YBZFOE(&4FE68fAU_)]9fVC4J)
7W2.D(f:g2ZPA]7Ta&C_/ZfZf[Q4Q]AME/[8FY)Fbd+IZ&ABGgD[#=_2cEJ<W_ZB
FVHGD5#U-KNS.Yf0.4f6.bZW4,-d=7P\X5e.RbFIWXXFW7_?HR(7#,</T+145F-7
+gf]#CDN1OGJR,U1/=Z[e?C\J=?^+I&G2&W[#Qd1DCCB@8U49W/PDPMcb]2KJBI0
/LZ1X3M[O1(?_/[W3SX7.3X9]BJ:&LePR3&::)<\,.A?PBf2(TNI#_Fb1TJYKGb2
EI7)=QVWQQWb-Z-](e^EX(gVdMNAbV?T[J9(A(/Wg-PH/1MM)H0@&ce&6]GH/_b-
)+W^G9S,#P[]GaN1:QR85VfFWM:gcPPg38J,@2\4H-H<Y<UUTMdO#H^OJ8=ZZT0<
GJ-7V,U1f&W;Mf,?/BdLSD=>,N^/K+U[OH,U5UU&3IH:fUUBg^^(\;AIV&:,9d\=
>L#/9O[[>a>M>0LTOHR;/T>&4/:>1S>\H6,L0)B0a1:19XS@V]CZU?_UeDOUVG8>
Vb93C?K4Rd4&U677[Y)[0[KVW^=P8b2;?IPLeEW@cS?+QN^)_;0Cc?ZTC3_DZcZf
S7J,)0HB\;\O.+e5.]R]?4JSUcKIL:e5F74\3?>BBE<5W6V<D1PK)0;3&Fe_DURH
U3^7-+UP+)53YKR]+5W0K,X8X^DeS8L8J_DA45JDOKV.D.1Ogg=P,DYWVe6d32Ng
6DNF53b5,T#:BY_cCEC=<XK9?IX#GWHR>J-5+()fQW8-_OSHb7VR1AF.YN4I^KLM
;1_[\d0?I7SDD#&+g.I6V\OL9Y;>7S.DVXa.MMT\Z.=<J)dg]J@<U,edNKG9H:EN
@6MK<eL(9=Z;M5deEB]AR7J=1g:7,,Gc/N^F[G3EYB&K+_B\eD0N]G.<XLQH43ZX
=R(=:A_Y=Z?QDP:G?X454#?-Ba\/8/+ZP=CL,Y;TB^1STeNaGLJQU.AEWHg-&Ife
fd:#,Q0=7^U^<Yd<(c:<K^-G,_YW-(D>S?XM6WGHM]4M,FFE4?O#0^R:0a1T=B6[
7A:6^CS#e[8::O<BLLR@e+B>6O#QH/M8J3D3H<+a:R<L&cZ-IIb(cO#/a0eQ4eN\
ZR<:f9RK;Rd>^79:e,NBE^O&#_SD9B;J0IX<,6M?SP9X^:.gQ+2&Pd)RI327N_0e
@YWP3-TF)XI&JR;=]3T&?]a1Rg2:HE=#YT,W9Z)C,e(2,6?(.VbaO.=(Je;O5f(;
I=L+K(#+GIN&W]a,FRS\7Z57ZKL6RV(-FZbYa4RU0_#L89eH3^R_Y(HGC;4[Cd<U
E8ZHg]T<^]XVST3VSc#ZC\786RKD(5-VRT-NYTH<3b-GG@@GM<8:P79KfO,f)gYK
.,gCT7\HY_RR?cU&RBDLX@?,4d>e;DgdOZ\EN>8Wa2LdO]6-=_5EM.E(].8IDgWE
a,E(Cc]YFLK)]J-:Q2JN>0W6C9d0E;.gGaeI7/-5.d3VYWH-^fF^N(_8[O^,VI(e
>,LR]WU<XQS?LaRc?P4EU_R_=gfI[VH8,OH0+]?WFC?(2#=;X04ZaX0U\CJ_1V_^
>bOeI(4EDa/g1Af@FCF6V>BC;6b1fAZ)V<A0eH7c6TC4ARYe+eBGNS:,-^X1ed?f
65<1J=)J\4&SAU7RZWa(DWWS_51:fcUPEG[1\[;D&Le,B(86Dbg;U1B7d^T:=0VQ
b].]KgCgI.)c&JP&?S,P[<.;3PF]F-QX4F0KVa#GH_A]gP+15)XL/2/[[AHb2RBR
OYW;88>DGGd:/ASJIfW.NE+)4D;>S15X13\\,KMfcQ/ESQ]Za5\V;FY;#-Q<4L.Z
2E&1Dd+WS;A#\[1SO[1dY<G7d9/G-7P(/0S^BfFA8CB<4dg)^.YRFDW\YfA@2O-P
FbLYegLFIN.(,GY14)61e4KR-dG(H-)7N.?fcVcKFBV5TZ0Z,Jg-]_D<aAII_O?;
BLFS:NC&G#)I^S;g1Q<]GOTcZDR]KcHK1SC75R/5SdIbbIWO8/cGYHU_RGcX(c@O
&=&#+=AQ>WaI.J>O2PX52CH4E.f)^DgP]cGBZ<caFaWR.;P<,@Q[Edf4RdK>8_6B
1cAe,?2/f,X^.E+^;&;I3ULd;>S037)9b<D+Y?:G,/8J0gDHCf/9AYG5(4Zg@CWT
gOJe_;O/7?V^P+OO=790B3R=?WN:Yfe>KV4RDF@/&3--4IG4CcGcZ#34)MX6Pc@Y
0eXKGaB_Q^+ee,N\^-d1aA#NAEO-U)adF5O&AWRgU5&cdTCSW#B(\f+9IH25U:eB
>F-Z)C)>;bM,2GD:/O/1G5)TN(Uf>8A+8[7HYcF45-5aGXc=.Y,2.4ZfMeNQUb[<
6EA4O4+f=Qg4FYFdU-#5LZ^>FD7aLK.L7g[#fQEF)cU^=c:I;Z7FQNAYAS+>>?OD
+=Y<&).9#]VO]Ub0X8VRg2]cA;0A;@);0-6;D)A9<G^WL/@<KIZS?271SF)ZI_Q6
<UR_+W1TCX\I1KC_:9QI?cab/(0(<@Sc(@1H8.3I5,9/,_,M[;4:Lf@;a/8QF4.c
E>;Q-KTT+5.@QfJDFVB9T]933Jb>=T.XB@L@?9O@S+aIUFI.S,-:NNI<K<-,bIP#
57QCO4_gWT:W\2MKdaKC86d7=0MP,R#VSDP>:99RVOYZ8eJD@8EbgR1RFK[>Rb^(
<Uc:+./G]:AT(Pa@dRFH3(YAb:N>c(WD7C]aL/5,d8ROW&?.]cBI-^Fgc#Z,7d/>
f@OfA4Q+U/1\U,bd]4-#[eB:=UE;N@>Nf:M+YCK<SbK+RJ5(ab^9LMdM[#F;+c14
>37c?0T[DJEcC6B<R-C<>5W_K,;\bC+&TTQg6,&H:1b??_EA<LW#Pe4IaX]Hd@W+
J(MBe6HYO:gQTc#2a]4J0-M\EF-JFIE<_]?HC+fOJQZLV#O;0Z^e_1_&g&;e-[dJ
cC(g5XJM)R7eY&cH.M1^85W1HL_Y]Q[@-UVINWJ=J.A/b/f;2C(.A^Ig1S0:@=7;
DO7LgYa-V?J7UT7dbaKg/dP:EbGVOc7Qd)4?R\?d/@2G]1DK(MR=&MV-HJKfFfV3
M#_A66(5K<X_<1d^6D8GeVeRV)Ta^9>B;PH<^,;2)beZE0dB4QQ(Y]5(L0.V[dJb
/FHa@L^KIW(YV2(gO\H?/AKGf5gMMbH=\6S#F^?e4aCLa1?@?TY.J;F\g/B67R8.
G\AI-X/LZdOH.PK&DF@1\PGC.PUP-DGb?NFF9C,De.547Dd?>0O2c@?])-^Z.0TE
egW_(7AW]S7BD9gYX00O&&-@\K=]<f5?ee<fHKT6D2Ya>C]g879-4,K4<5I_95&W
_&W#c>M)4GQMeRT<40bL\dKCc+D/FIJ@eDWB/98fY/UQX)ZdO._EKEEVFR[:]6-e
YG@P]afU@;)UTD/4U=Q2KGV]2Fa3\\V.TZZXP.ddSecD/:dIX(&MNK]YGR,];_EC
&]J<G9baeJQ,V<W;)?O6PW=L/I<8cc1U8)IN:04#.f4b#1b5d:0+V1E97?XV>-cU
Q&2>,2O5HSQg+,A,OJ^VAXP^GDG&EbPcggPd6+&-/G]0THG+]1<[[dT=[K)PC-fJ
e?HZ9A/+&.PeL;YcK19DWMU+TOPH3YK#]B51:Z\fG7@L/8cOaa:gaP.X]Xe\1M\K
W(UYa<cefV5+9NBQHGV0W6&5<.R_MHAF0HJd5Gb_#6Z6Q<9>G2ScHLI\b0MW5/B7
@)\X5e^;#Kf+2CbY]dQQPJJ+6LF>B,7a+Wd+WNMV>:;5c52[:,Fc06.L@[c;C,<&
Mc;XZG^YR>5ZB=NH&:[<P>2.A>H5d3aLf3(Ha2b_6IV7aM/e/-QWHcWJTRP+1FgN
A.6J1J5@,S;AG\Fbc9^5YZ9ZDK2f19-c^F:.;].HGV@:eKS3L,^dXTJN[V7HJEH2
O3^6;WfGVS;NMf9E)YHKYfTV0MB\;1R_?\5?WR>Z40SO2ET9^&8>]\9gPE:KLCHW
7Xb,(-RDT?gQI#(;Y]7CM7-MXUFFcG^fOHQd.O5;aQAX2aV0AY92K[R[B1U;DJNg
aU(gC@5J728:N3U5#_3<]1#Q1AUJ:NT:X^FK,1+[.10D-)9DB;#4Q#J7;+9b/6^R
f0c[\B=S5@?K#-8B\bgEScMQbR\3>4J^4.KA5]SP/RbddYZ4/[,CVUB@/8N]^P+<
bc_1#<VI;CQ/9R/WOVT-\^+U9H9K(DS+8K)AN)3XEXd2=TIQ;cW]P??+&/<=3C&X
D0_)\b?@afXKXe/c/3J-98/:<bPL#HW/?(BG:b9<=L3^33M1FY,;5TK,15A1XYYK
(Aa;R1/SfaK1(B3[BVE?C@=:F15cV9<J>N4T&7&/\8,1D/b]CHRg6QDf>]-M<c&2
W1a(E:dG<4Z&Fc^EE?(V4;&U5e.)XR[-c#Pd8SHCKdMd7aT^Ea3:7/(gI_5E27=K
Obg;f2a&+P357T==;_85U/\4R),555c1-@[@Cb-6GK+ZE4N^9<NRESG:]_@<EE5@
A,FMfY;4SXgE?L6.ZK2N1BDK<Je?/;@_KC@dR]T-Ldd&=/0P4/V81_aR43M^-3\5
QO9YPR;#(1Ze5/LXgbU_RKN3M/Z^VT(&_LQWN#^?U>W(Q6.RPYMcA3748V9ML;C(
(G;4\P^9S+FYX-CN?aD_&e=YTb?QcJUY6P]\dK;K7.R;>a7ODY^4Uad@7:?LG.)4
_Ke?[<ac4I@_JMTc(6+GgA3dWd^/D>\XS&dKOBV2g^J)6d+<7D1O5R)4J=AX1OG&
9_]GX-39WJD3WH]FaN]aPD5I;/X8/@^9AXVdfcDIW=1<28PcU?^OBFFB^U>E/4GN
)S(.P-D9DTUCf0#IVaK86N[ODM0_e?83F2=#_RQ0dA=DA^8g@:D78Yb2V6HA;0XM
D6&D0-+0RUUe4_A:8F2b9G6DAWJge2e6=@^347)\F)3SCM/?>W0U&>Z4g@E75^I^
4:](36/WaH101R+&V^.I<6:R;+.,YO,Zc4J]:Q[4F_>dU2);2;,#5W2/.>3HMC4T
-f\A:=\<(-]_1NU3HW1M]M/g5H,\+JX0VZ:A954aa>Y#E:.WYDdcb8\A0JcO0<.b
,_d^VcRH]W:@aL[,+H/(/C]?e]?R8Kc-;gJ^@J\61N@85NX>4f0&Z(].Gc]3WM.B
@5AI[]FbKYEfd?J@8>_P<L5AM>]+gUg@K?/P:aU,YMY.<KWZ5ZJEgB3R^0LK]eO(
8dH46N\a2J[E+:=Td@+2D0.=FY6OUZ]M1+2P@BE.Y.g^EL1Q<;H@QeEP@(^75&1;
);T1H04\MH86=@):4;@CQQ<D&Q>;TT=ATU0T6[491GAA#D@@--KY#&_D?7g+L8dS
2<:-T1XEeMbW,C:4=M^.+])6e&>(H18eA8]?D&[GA/ZKA+6PGgMfFL+[/g/UQTa<
UL45JGN([[&V)W6HJT+S=d1V-USG[aEJ9_ST(5f5)9DE&(:AA#@K7),J,9KX&cX[
WU/NUCS\U7G>[0499#=HG5,:)I3J9XSXLSET.@_&:=;d=]f<A/R;2L:/W(&?M;8/
9G;:L8C1=WBbW4,=Uf>/]TN+?6PH)^#O9&5-_,4ESgZR)T.\0>Z-;R(#=D<@BK7U
LTY6_415O<8AecWRX4I<7cDf:@4IRc/VTM>NI=gJ3,@C[S<dX0cf;#O0,-VZF<:3
(HgGQX_\6JWB;8IE]b6cV\Z(6?LDQ44)9UfXT7LgGYJZTM>E\^N7;-HYTVHadHKA
5QVZJSJ&2GSMX(b6BFO8I(+_EcS@\X5-J?fC+1L7UD:K+(#Pcc@+LCXD)-VS]2,B
FF7JNGZ8RJ:N_+70>L\JNEW,_]eH:FGQ=F]OBBL66a5aT#g01TH]g3X\.JV[RK[d
#[/NF<:>C8FgQ?M9R\GbLI@C=DdBQ=V+3/3M+\5O1CW./UG(>YC0eOYaaRUB)+T\
f7;J+SZ;F?528.eT<ZOLBOE;8-I;&0SU9a6HGP^-I)=5dAA?A0MV=<+Z;MgPYM29
W=S4Q8.M/&XNP4,C=HZ[Y3\A:e&YU3F@g@K0O;1311#(fg;F:>e<5TMOHb8O]0-Q
5=WS69J12<LKfRP&BW)OR-->P&/O(WZ\L[d2b2+bCefZbX\EO6.SAZA_1V@B;OT1
Yd3&d7=&2<^5#)DSd<5X/;+I^3IKI;-=VRgSUYD>_aE+D</c?UbV54/5>/F.XX?8
:f&K>C2d7M/0]DUZ4d?LTfLT]GeZgM#8=CF>VT;F/eV4\=TfGK6(+YE3I/O,KG&8
2_S2VC)JP8P]5,&93@Hf0FEAI1<_eV52FA]]GP&eb74ccGES;AOdE)-aCffIf_W)
?e@^IOb]GaQ1XG2RV,_aDf:\4:2X7M>;N2<7]&FX>;^AN1aLF=P=e+6&IA83ae#&
F2,4?];+(:L-<I4XQPMe41gUMJAJb@3PN[8[;B[^X9VC=D#2NJ^^aB.SK2O-aIg5
5:GL2?eC1=G3CL[4BOVSRH=JcD3d5H[eT5(Y\^A]E22fC[0X_KD18]:#-DA?.Z>?
T4#3\K.A_3RWYS>-O\:0I=BAPZccV2JGAf\d;@/9#;\DIeP/Xb&M5:W\V8LaB8K\
2Z/Kf<C@>c\8Sa46T(.B+a;RgJ,=/9C2:1&:^+/a:VP^5a;NegID-5&A_MSLW7=U
JN(&:T5>)d3GQ+/a\\EI[C2G5[_\852OVgLMG_OX9,#YY=+C,L;&WSZMDF+L5/NS
FE3)CU?Ab/2>:G3RP-C8aEF:>UgdG5d.@EKYdRJY,PbEX-e,P&QT8>P>J1<TL0g_
QLb31@bE/g@W_ONYJS-GQKSFTa)(LG[G85dQXZAeLMR3Y9LIAa;P[KeP#42HJ:eX
&ZN,:^7dNW4[HeV3?QRZF@STN-)+2&(-^aKd^LI@??:IO>1J9J33gcH&B\eX75;Z
6AZDRH@P=^CdQ.7#>X22dAUCfAMBAY:NIKYS7>WHR3RV.Wb6,VMdcC]?F]L=f7\>
HS[UKE7P(Xf[O7_@<E61_?73UaQT57ea\,fTHFJ\B[f5>8d)Q.cM4&=7-#2^6S<R
Gf6)]=_U?;39).39,VUR]6VDE9_)9ETA;OFMcN+EeNfLWg7H+Q>UW1TVY32YaBX9
\ea;38fH]-O;PNV?_d1QdKZ<E?Vg3XM:,[ZFT6g,VaQ6,[[J&Gb&/FQ_4F6XOPZZ
e/Q4HY7W>=3K#FT(Sf(-,4KF3&HTM4X?+WM];Ng;2+:2O2FGUTZdeAJe<WY[:L@X
:bUY:C#:&8DCI3SNM8PY>AK/CRdC)Rd&^)3MLWJ#ec/2=a@TN534Q17Zb1T]GbaJ
?\2gFdR3HKLRHc;DBcI?XFO#Tcd:Z[RA(\faUdA#[J\QSgA@=CP_cAU<SG7-@+[1
T41/<4++2cK-HDgZ7)7fYR2JHa7JYEL2ecXSc/.e<]@d_;FC48AJd_ZVR]GXWcLK
OAB@Eb^KF&f3L?:5+CZ0LbN\E=GQMI]bU^_b&Y6]\5cJWe?S9[#./8NMC^-fUL1\
,#58F[LVVZPde3+=H#;.T<5N(ERbC-;d\c]Ub)QJFZcB3W\TXU?.aT#1aQE@_L0-
<S0[ME0#@(f-[<(VG+YNa8DfB1g-a8-MA]>=]=T5f&.c=1O&9b)4W2b5QT/eUG+^
#aOG.T>=5,I1a,A7&PR2UBK#XBU2_E(_5E>)G>0IG+/]FMRag-b1Mf+g++ga4LK+
V;;c^E6GE;6I5^N@bBI[.8<PI?,;5[,G4FQMB(_/=@/BM;<2YI)\4Q+fWJ];D2#\
Mf7<7ZU3^?PE58.30LKQ_;:Y?W=9UEaG;0^&cRYIG5685-KI]BET[/?0@c<Qb_#^
VU4/:>G/SHCNJIX5[-8>X)B_N8)C:L(d5c1_KK3Je7.2(IT_IdR8M@MO,e@8RFT9
aUYTH<fbY(;+Lb)c.EPTSV\Ec)D^76?#-6WDT)c54A?T9gbb,gg]TM-2c?@EeOQ8
IVgY<D\/]:TQZ>H&E-_UQK/[[>C5+97QB039O7S)fa8R470e&;0P;OKZ4T.Ace>;
I9&+W35OMb1,4-2G6)2UF^;:d\0GY/UNGSDG^96RDO?H8P-H[G9_ZS/E]H34MN@9
2ZVW7@3Bd<\M#[X648McFCH(;#)3cBIgO;SG@)81)Q<P.G:.f+SGe+=2R&3;8ZLI
@?#6F?3/QRL1E_#YJU;2U<XAE.NW+CKA[d).@5I;Y(&CI-+HP+;\@PM.M0<M+11W
VcC:L<\4J\RN#<NZ[I1,@ZBS;4H[V/RQO@HMdG-NcFQVA<bKE.PG&2eHa.UQ-?G2
&8eNG&<@-=NTWN,a6<Q@@Ba1VOW8bT@ZbaR6YK\&@RXKBD0bFUL<>Q4^^dE2d-]J
A=22,Q&3=M-M;C71#(bPJ]46.D[N,1Ze9#9U2>@A2@RLF^2YDKEWM+:VH7#+<[:;
)M\LR&B+EBT:-d+<dM96@YHV-X(baSP+2DSEH]-GP,1E,g;.HVR(dSR1=dg?^[)e
J[7&Q1HAPD1Z6HA:F4-;^.^dE1Hd?0WKBQL#b=I\1W^^VVR9WRg<&\LNW1D^N7Ng
P.0VAEV.=eV48LC;)1&=VV\g_RgI+GF?e5<G:Y]UA+ZC(d<_ZV&E^aUC3GP]6,6(
Y[7)[J61fYBYa>-LV)6V0^C=L-:SUddW_X2:HO9GcSf/R+C=6UN?ZN6:g+eQ)??F
[B3F:??ga+OX=9]Y-+H?/Vb;@GccBUKeO?0,/4YF)Ag_g0Sa)7JQY#.MOGLWWX37
VBa9WSDXU0P&7A^AFcI+5Wc.>;7@NSS=6LZb<_J+#5#XL0_DeLD?Q6d91&/A&D(c
NGWXf;HCO7J\\c8+>4dU2Q^E6C,+bR3XU2FOPQ15M@e)4eCEN)XV.02aR\S6D<dH
=JXL>>CN9=U1GH44GQHS@R12>7]]gDI8HG^Y_U[<9_Rb\./HKA_U^#aU5?HV9-(e
b<9RHEP7R91b]\?E7&E\CPU\ENV1?\eLKNC[cV^CJcL2g_A@A.eF^^IB.cRBId]+
S.(3WfM(F(g:e:NLGS[[bfW:W^W95g88?e6&,VgPUEFI0:e(:)AK?4ZXN(AO4Q1C
&3:f8AFW62Q/)^g0bP?Ge7;5NDBFMQUXO#aS3Ad+R4@O.@]?DA[Q[DS8:K?Ud;(>
+[I2fJ1:gc0>^&H3N@G=D5^4F3NgcE-<<I(A/W@_RX_V9WgI^<NS50/T]RV1&1FM
KM;#a[4DO;7AaB];/3aNcbIB\.Aa/AH/DL+c-cC7NN1I0Qe[?0WB]HWUDMb1PEQW
I[J@>1@+R4HCOC-T8?.VbAc#IES),Y4[=V>CP[,9,278HfL)KS5Y\YX173J+C(3Z
>]46BI3^#>+)RbgJ#W1dYXOMAJD[1O3+_,6AIFAAFD-WVT:,N+-;;7UcKdg-.f+J
T\N&0PSf.O\&I:8JYa=S5#7B6P(:^^A_WQUSF,aQ-S.N3VYZGV2ID)[G61a+;?c]
T9HE853c/Ag(<HWf62PbFUQf:O(V\SLc/[aE_0YDAc58)5.:D<UZ;3gC\F:]_XZ3
?[Y4_4=L;-Z<TN-O3\TMSTOWG)/3F4?^Dg[S.R=#MR-03/\)aBO5Za]9^=bW+0V#
C@XeM?C/dfX6:ILZ&MfLMc/<ga@c57^255PRY6U0-PMH\W1FM^(@5T4&8LL+S30X
OGE3F+Nc8fU4EK+Va(?;&4I;.^3;46J]c4#(Wd?>N:S2/--.ObOF3;]O3JLG557F
+HSSAY?&3).7->/9K;+&\A9IHGeV;e.+-_;=[E4NcIWR\dA7VPWd]75Y;^MMd>ER
T0FN/G3.2II>/-dNN_bBBWU7U5/-6f?9aZb_[AC.=W447X<T&Lg=RY/1A1Q(+2HT
/OA9#=P(AQ5RdgVfDf:Y5@:DY34&#-;I?B.?=R1Z3[e3X[?C&R9.]e&MDC+3>I^Z
JX7F&76)IEd2N=^5XTR5#:TXNUU[:Y7-JC)W&:Dad):BB7#LSUXDd\L#M=bR#3XA
^/)(#H15,WQG\]5\),GG)&,d4:KP]<0gd2IJ?bS47JTWE@=Z+ALaIX#J3#2Zg]#E
VDHe[PTX4b05X\LAUT5(NQ9fSLXdZb19F,Y,DPY_ZR9ad67Z]=CCHMe8F;GW>SB1
L_4a:Z6N_H5]CWNPJWfY(M>Cc/COZE:MW__.10B@Z_fF^]#<.\W>9\Z@@eXG(NN-
NGWOY3aMDfd)g7\ZA6DXB1XD9f7a/,7YNBD?\IL>Z\#@6cbFYc/NfJ?=+fXG)=\S
66Re+X4JXTZ.@7f4P(aYUTSB8BfdbcQ(]D(+6#C8WVHS(?HZec^(8F2VXD(a)WM+
ZBgQ^+_0-:RfTdd,E>UX/0,?+4NZBdE/3]c3(eEQG&]Fb6J.Z:3SG[/>TOIOE[Z3
@G5W+=F761TS+&O69YgG_5\a+TFDHDG=(20b?V<HKDBBa3)[bRXZ37a)H][X\3P[
OcXgD[L#_IQ-:Pa65=G6S::M5>4a;AM]B=>:ETHf@324d^DXZ^/5FR/KC)K[A^Fe
8[TP2aCZ)GEI,gff_X/0^<^J)1<>)G91[N\&VTXQT>D.\ZX>5bd.Ne0XGAK+ERZ@
Cb@M2MOLHKE2AC;R.Ae\,:)dA\>g#BfGY[2KHOJ4C+<.U_]E-(aR=bFQe7a0;:Qd
a:@MW@fXE@<)1<&:Z&7=DfO6ICE;dNS=IcC5GCgF?#b-f?(\dZ,FC]L>\?ZBKX)O
KdLM<Y(6K)5GNIB,^dXW@Z5M_JaaKaK04KL</WWBT6L>gEGEcfJXD@9\^T2EZH?4
:c;G@KdF4/,MA8,WXYYM/KJ<D0T0eLRFYSSHLgJ^NC#6V3EL\SLHcd[XdTBf:B4E
4Q6[AT<IQ1=2V:c;UJQB1(Y3QY0TXA67]3LO8QIS():F^8g77&^]T_9P3].+\J]V
Qf8_P]S1UU85N<#.0T9gf1a4AF0_+](-OL+;.Ia.2f7[/R/IMfa/O^ZOXY]\@YL.
C;[;Sc]J_K]+Eaa]OOO-),C-R)R:NUgM6IV&)TF\GQ7=De[-5&UJQa@6GeKJ+c9Q
6d<4DA+-].1T_YfY\)eRHAL/T8aeNZZ#&<8[>VQ#1Ab3&2eA1)BFgD9NdL#77YV/
MEb809=(P)I/T6@a(MQg+.0;RbH=9?I@D7\];bA5<@TH[J8Da=+IZK_(,eG#?L;g
L._@;f_SQ40eb]Z<T7&=fF+JV3eNX4_TG>GaB??.X=f9>)M#AL4VSXN\;K8;+;9\
DO[WWG,L+H8:5<VHN]VV31FER5+O5D(-g3gGe(:R2M0:&M0)ZU@/NS7SLNIP.P@@
VeE3b63a:0]M.75\5XUR4FR/4[ZaXcKC;f/RL6GTFd-A./O(b+H15O]_\Of6;Mg(
<4>+TJO_(/K8^9-Y<T5T7,?;6UO)gQQe/gZ-#3,RK7]D;<D@[.I/3[3)b&VHA>b,
<Cd>MeE3T0,[W&\;QHe--D@Wc8fcVK9CKDb(UedYaP;N5^T2UBe6OcJc0853:,@6
#1S(&D^<[96Ec_).K3?a((9#KGAB#&)__M8^:c&8#=KU@J^QVQ^?#OOJZLNS.<,G
Y2Ka-_ZUWI3;Y/3<H?\?:e7eV(VRXJGM[X4TX-9W=BbN:Ma\47Ob]IAPA#).8e6]
ULd^aB]Q9T:R4\EfbDIN>MA=PR/N_B]R3#\f8L,Y?,UYBLC@Z]K&=C:LT&SC)=8?
_\V(EK?d2;FD_/>-dUNJL12>fa]WTL-Og<2??XS=c_6OF4MdS4>Rc#G(0<TMLSQ-
C\E,=JQ:2V-8DZAK2Y12g5KK;X(47Q;R[QNUHA#[f1;50E=C5.<.NY\?@;aR[]+.
UNfIJA-bS2UeGBDfB?=/[?ZS<E_T9.AQgI1.(+@Y>V^M:^ed<bHGeL7S#E8[1A45
gN_.6A)Wfd=gY+c]aU;9d]F=,GJRLc&-f51GSN/2ZdH(V:A3N-;:JD2S3,28cX2c
b]bcQ-?]/:5U3=b6LeeK&MG68J?775++)ccA+84fZR14bJN]ZPbH[G8fC<(Ub8aE
/d/DC^5bA6\<95.IaW26c?<25#^+--A5eP[V;N8^\@_2N)Q5[fE_;5@;<./,+[XC
/YN[=#c7859g+8W6gTPcQIH=7[8c,5FJW,eW94-@4TCdIN;@ffU0@<b+bTd1c9;9
PA=#TNB5HL[9P+YL=+:>_G+WY+=G;JfTWe/@#0SeQXS)2+#&3D,eU#5KMX7DNPO(
)I>(OQ@HY.C2,12-GZR]BX2_(>R[.KFD>?5(IOPcRQRZJKZ2Y(+^B7:9d2WJf9KS
P;AI[UKP.X(UXN(TdDd+M&QN1QU:&22S;c.CFeV;L(X++;gDZ1b4Ac;c^SE_>0WB
^?PQe&9F:-35-S-[dIF=\B5K:-G1\B=DJ)-)N=(K&I\^8)ZG39\T>_D<Y&>M3B?a
KfF:7G.FUZ3\,5:bLaXP/MG0;e]@WfEXgOX>-[23)(]V9edO=CD_43P\ccOI:=Q]
c3CPR\.]1&:2:/6AQcT2U21XC,5+Bf7bQ-Cg>VRGIc8NQF-3Z^#OM>BdgW.<^Q\9
I?7]+INXZS_Ea6FK:ZbT-=?&T+VGQ9Uf&Ee^XR8gC@eGegAB6Y)NK;K[6+DE+7Fd
-:^,[SO?B^_5TE#_I.1eO,#0J0ON;(cdPB4VBJ3?^Sd8-aG^^07A>a\GR:GXXFaJ
79?a)e7gS3eKa_G.1Z^e9)4#<J2F@UD5BH2+#>IK^6=M06\-OEZB05bc83e/N#[9
DBTYG\EMZ3gM9X,;F^[RJ-0b]S7L8,J8Cb5^HDM]T5+BV]8-c(,N4)AG>J[K>KJ=
IX)<Ec0f+d9D58c0OgPE3f.?X(+&LFEBI8:ZdF&\PPP+=MdL^48C0I-O#DZ88?T9
V)F^B=C6#^1(0&)9ITF37O4Q[R5cdHGAC4bH8LYO0<+aMFAEDeCXO&[fHWP<a@W>
d@26d.SUS&F7]NK7A(VTC1>^2J<:CMKL0LYN_JeI,.-=58U49ISQ^>2We)]Q/U4^
C_g9Gb+/+&/8QGM8AUD(cUHa0QJfYWL:#92.BSgR,g0I/EOLE:a)OMCPcM3?[A<>
#,SJOQN@I7K[bcdbHdb9?.eE4[4(T=TUV@>NA?N)+5L4OX)PMBZ+@V=)H).Z7,bH
+#P_3BP+<#I2._E[WTe3@3LO]72.;LX6,HZ_f&QWY^PVI<N_[KMR&AR<F_<CGW9E
]>/R0+g]_@8Cd_G780b@CTAB?g<H305V/9E27N\C<5Y.>a<BEJ)RcUWOPY@3aF]^
5=e<]@+aIZaEFI9A>O-.KK=?cJD-;#1/#N39.-^<[N\cY;Q4L6C@HfWU35@DSMX[
A)6?T]JU(Y<2;b6;f)W#+-/A0T,3W1F,b<[L?=5b7_-5]#-/>6K>)S2O-N;LR/CL
gOT7<5Z\c_cW<5e>JH,f8c3KLa4EDBB1C2fB7W>:1WX>Z4.-4HF\Y47CW[OH.H1,
)aRZA?=,V],.&2X]Ze55,ga\ceFcTcN,K1_bYWN353?f@B?><B52]dKO<@aN.7KL
,,Xg^R]9Z[1IY.&.XI0@4ROQO:_2GK1(_F\J3&SfOM.)CLZ4XDKV\dR908I3.E@c
RNc?QSg)3F<6/VO#ef+LGd\9_)6=)g0/N2He4,IB99TOId2Y98NIb\V2.7XD7Paf
CfTWL5E+gDCRJaaN#G8-/=-@?C[&+Z4UWAR[AKASD0YPdG[01.^/TF5>&L2(geZg
Ob]NVga\aI3YeAIRe((K#_K1O8bI()977TZe^2a1)^]Z8f[:-1(1OQT,\G_Z9L13
13e\=C6KJa].V2-<954D#8_Q_T[L[2XY3WFdZ#XZ5WX5+L/Q8#?UYf5AJ3](VR^c
eF3GZ[/e9OeaZa35FH+.A0K:[CM]:QVdA,ST^5Y(?f/62_4fA@C,X&4W4(I_D6=J
[YeXYA-TgEYM)A)WG)+7S[QUc4MWa_A4;[SBQ]+<CJf]82_RF],#HU@2QP)W^(#V
ZWGY;MRV^+:3LTeY5^?XJ-7Q3?D>:&)]T/4BO1aF+;K<>be,CacU:P\c.c&=@.?#
BI[CVUL.J9(\^CdC2@EcgC4Re[Q3eMd+;:7U32+,d&3BKS,Jg?f;6Qgc7cR2O3#X
Y1JY?.#fc-G.[9UN>7cVce?F1)Kc&?+JNLM3HB-4Z+OFE:0L1U<0X/dCI6HHK.f1
SP]^(b9U27XM,VbTYUNL=M>JW_BH>fVd2:)8([O-_]_BfDe70a+ObW-L,V1aE\>]
-R;+(/98L:QRRG:cV+cQ\J,J\OG_<8H]SG;V?Y)U)Pg9U.CSI7YM,,)V(4/^5Kfe
]_F?5c\YPa.Y)+7b)>cSXT)=Kf<6],E_D=)=>3\T5[JOb88@20(<0B>1H.d_M?6+
2SS.X4+;0M9U#O?<HEYT:dI\;B@Ae+gG1ZL)<6U>.6P3-;c:0ZHCR[01.F1gaX3H
g-c2TFI2BF3?-QV^ZG()dR?5-O_,<c(HRA&S1EbY,ECUEMbSO;1N86B+<LMJ7c9d
XDM:KW\23:D8(<e),e=F;X3eEeCeRNU5AIVe)I(G=5XIIcAX3g-\WYK_BWOXBW>T
=^E\\[aNg.XE5XTO7A.\[@/;.\3,@LP1-_,<#;@TFJa\[?O,ICBJG+PaIJc96[C9
2?A#;EKF5/.>0?=^NNTI).(FDK0WTbH382X&L)#_9\SH2UE&AB0QY8>6.^,Rc7K;
1=5)6OD,BJW+7F6I]:Ybd5&fF0Z-JV_>H3c/TUG<C:Cc_BTW^\EJCcKHdUB:Ob,F
7Z\^HPf(:?.&8_Af@fcCU#(R0^M=K;0dPLc:8cTB(J_W.1NbK1=2M.8f3S+G/>ZP
^7NM?YfN2:I@C(&0QH2IJVOJ,YQ)1:7fIg/>N<._V++g_6;8A?GENg<8,K6.:SLG
cCXcQ/C/9UBYY[=:Ve;-\f).,\F8<4K8=_=3??G<c<E:b220H]\aO-]Y?HR\?]Pd
XM?b7<a14JPI>>=(ZY_G_N&Oe@FeT1/W\dF)AM^e@Q.M;,ST7e[7FO3fc_CQQ1La
g8B.g(KSEV3G^FDPA0?3#-#B5Z]6>_6RO,HgDeF=K8)5.5M8^OV/GX1#^X@7/<-]
ZD8+<?.I-R>,c[NBXTae=&T.;L1(Dd+6c5K.8\>N,9.VS&KMS+MFXEcZ[P6#XMa8
Z:TMG7.QLRPCSB0/H#2S\=-a]TWXT-_,?Sb\W\@Ua)GIQCQUO=,B?9VPWI7SS[0c
+YNgbHG7Z3YIe^Dca7NTPGW-+K)6a<1X2,KKdD5Pa^O+#<([<BC]NR7/)2^#NDKB
X@^._&-Z,15&S46>^WfO7E2[LUO>Jg8e0fJHJ0O)Z1&#dSAead+T/;[@=J<#LDbU
CGURP:A(7E7@4H^B;32GUEV:4]C5Y5]^4N/>,R+D(fg\,eQ^&/4-c;/X]d]2cS]N
I&>I1R2UI872^I=b?RYHf?c^\/(69=:DH,(CRLXN028+bE5,-OUbI2Q23^?9V,4f
MK(#G2XfOXReE0bKMDDQ0Z^=MC>\KR999@DTcUC:E9/8L2),GU4bR@#IA.RdJ3N@
01UJMF@]6<]63b\NO+IWK(&A??ST:&f66I9g,BOH/dW<D,gH,L@6e6&2AXN2QD2Y
?&0/8/f50f-?Z9>58CGJ&URAfB.4d@<+DKO6J@>3,7)FdM7-EaFESR>-ZZTKA>Z3
b[&Hg0P,BH(gbOV_0JAJ,PaGE0\1dQFe#FW2)]_=G6MUaANZ)(NQC(#fAdcKGP[:
=&,L\L8gJ\=6YK#eI72GYg@CgKG7Vd;&)Y;fN2WL4L#ae-B0[FQ3./<C+<gWK#CK
5cacO?60E#0]?04)5W;_0EZbKbdVeV./I9beKCRS[S]UYXHEeQ,UK\:K(GeA:I7K
UA5]\RWX61&R+XPGW;W<Y40+99T6dYR6a?5.WO.2e09GG<&C#)/TdO#fTf)Y/2J6
3X^K?MZ]JJ5WWg=M)=V(3<]KR(#O5RbNUg>7ANU1OG+II0:+/9W^&b5<?T\P]FDd
1:#agCR7MI\d.R:ZK\_;2.Tf[@+(MVQbC3W-b8gGAFS,3R_)[7&+]N,f5\99E+AA
=>8P\O]XTC(UEF&<3YE4MA1?7VS?8g@aUJ9&5YNT<7K,WRIB.3gd<(\-9KSd^0,D
UA:X6MFa^8KGK#]a]U,:]aPG@?HFF0O<9b3(Cb[8#[?5\08dGI]+bD<:Q_Z-bI-^
a6PH2aH;^I_fabfCCM>XA+\\aSO7D:cJMe;f+-Rf_F@BC(\E?-fRPIda&T=GM,P/
d3De>#>EOWDADC+97A+4^Q;H[gIK@T6_)I2U@<>=WHQdH3bb#ddB,7P5^1&JBa/_
9@@3NG&02D)U,?[gc/RL_fE<Vdcb.J9[7,Z]-WE;81HM/?1@F9-Q+>;QY+YTH)M1
fCYT2XYUBdf@J(J,;Z+6J]CCY_g^\>7JS(9=NMecKbET.dB0Z>Z1?d;a)13b>_AN
129I2@SNHWE;,J<a<G_KM=RI0aUf7H@6QUS?.-f/F?(bLXg+WCJ8IX;BEC_^dVNf
WZO4c)3^gP?cZK+T3M\VAG[<[Y+S+8;Af0Z8eg[8QF<DA7BJHK&183MJ6g-e+ULB
&Q+S^Q#DX)-0QA<Q?HN=@:#AUL>A-=[;&8=L:J9Z?F<g:L1bWSU_aFdC<+#9XQBN
N)?UZ^ALG1-,FOW3H7D)2gL.6f#=PKgXAS\.>,X3DbPKeb6#V#C[KdFBJ7KF7<0K
3G:c:T5Dc=9^.:I]K\>L4(2_,bS2b<fF,4WX#6RZ@fO,2R=Z#e<8WRMDBZZEU4_Z
.E[0FZ/YYWMSPPdZCXMMQBP=8,0+I1/NAE\>(c#-KOX]URTT8bW_a1>O^8OUeCEc
NG9?)F&S[GZ6fXM_&O0;W[0W]6[\BA.R1dH=UFKEQ\\]26#)IZ,4B+TBF=d85-.c
T,Fa^9V.[V05[d-3J8X70.g;=:.(J^,LUW_)ZY/bLE.4a4fE(1)3K@(9IE(LD=\>
5eDd+3?^MEC6VK2Bda6L4>P4\fL>YM/Cc865?2SKK.N/JVHW^\2U)DK\GOMDY<.e
S/V5KJKaTW<J#@0EF&e/C]8ALLH5MC=2P)-fZ?cE8?XZfK##JDCJ)+_XR29FM,2a
>5T]1;[g>fA3Yc-XL,7)W+VK0F4d<EXP.8^]VXbS-OM9],\#d&8Q,O.@b^TeIQKC
ef+H2LL7CA9_ZgE4X3eI?cf8<;WN?^E,5NRA7=IO?TS\M1ED?SJ[Cd+++F;1;[1Z
#U:>+2IgM7dAR#LKdf><QQ\B\BU\U#-3.aFHO-Y0C1)V<5PW3:RT[F.Va)KO;G?&
\^^7?C9M0GgbB#Id.8\,d3GP8<ONQ-V-0>TG3WFLfcg?<4f[58P?-dUU7fFCS^Lc
7S8,^e;YTY#HT9H2YgZP?KRcK:2@3^QJUQfb#97UX&(fGA394,56OaA6?-5Lg=P4
9Pe16E,>H_cF083P,@GU4+fS#aK>JQ(VJ6.eO1V=LO&LQ4\253J#Xg/DSEgS;bB^
U9T-ZU:S=U6L-V+)fcXKD;e_^+691UCc/S<^N<NR@?=7/4bWf&Q;ZQcK#DG=:1fg
3HEKV6cGSH?aC=CWbRN[e(V25PB2+)VPVHAC9R9C3A]##<S[JaHbW@eSaZC@F>E\
9\:]>+YV@cP?Q81>5?B7>cTffVVaUCaX4U/IA>PHB#\aM,8dNJZeMd?J8,6/8+UD
LYUKCCZ0=SZ1b6ZH@[D+;PV;+BQ7+SF]J(727AX(DD?9SG,IRH96&+XRWHFgAfSM
3aZB6eQBc&E->?g.GGceCZB];_7Y,C[#FZS>)NV=/?QgK)/Z0TX/:<@C-&9gD-Ne
\3XC3bX7[T,-+$
`endprotected
