`define CYCLE_TIME 5.5
`define SEED_NUMBER 19384566
`define PATTERN_NUMBER 1000
`define DEBUG_MODE 0

`include "../00_TESTBED/pseudo_DRAM.v"

module PATTERN(
  // Output Signals
  output reg clk, rst_n, in_valid,
  output reg [3:0] in_pic_no,
  output reg in_mode,
  output reg [1:0] in_ratio_mode,
  // Input Signals
  input out_valid,
  input [7:0] out_data
);
//================================================================
// Clock
//================================================================
real CYCLE = `CYCLE_TIME;
always #(CYCLE/2.0) clk = ~clk;
//================================================================
// Declaration
//================================================================

integer SEED;
integer pat_count;
integer i, j, k;
integer exe_latency, total_latency;
integer f_debug, f_dram;

reg [7:0] DRAM_r [0:196607];
reg [7:0] DRAM [0:15][0:2][0:31][0:31];

reg [3:0] test_pic_no;
reg test_mode;
reg [1:0] test_ratio_mode;

reg [7:0] pic [0:2][0:31][0:31];
// Auto Focus
integer contrast2, contrast4, contrast6;
// Auto Exposure
reg [7:0] gray_pic [0:31][0:31];
integer expos_sum;

reg [7:0] golden_out;
reg [7:0] rec_out;
reg check;
//================================================================
// Main flow
//================================================================
initial begin
  read_DRAM_task;
  reset_task;
  for(pat_count = 0; pat_count < `PATTERN_NUMBER; pat_count = pat_count + 1) begin
    input_task;
    ans_gen_task;
    wait_task;
    check_task;
  end
  YOU_PASS_task;
end

always @(negedge clk) begin
  if(out_valid === 1'b0 && out_data !== 8'd0) begin : OUT_RESET_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("      Output must be 0 when out_valid is low      ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
  if(in_valid === 1'b1 && out_valid === 1'b1) begin : OVERLAP_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("   in_valid and out_valid cannot be high at once  ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
end
//================================================================
// Task
//================================================================
task read_DRAM_task;
  $readmemh(`d_DRAM_p_r, DRAM_r);
  foreach(DRAM[i, j, k, l])
    DRAM[i][j][k][l] = DRAM_r[(i * 3 * 32 * 32) + (j * 32 * 32) + (k * 32) + l + 32'h10000];
endtask

task reset_task;
  SEED = `SEED_NUMBER;
  rst_n = 1'b1;
  in_valid = 1'b0;
  in_pic_no = 'dx; in_mode = 'dx; in_ratio_mode = 'dx;

  total_latency = 0;

  force clk = 'b0;
  #(CYCLE * ($random(SEED) % 'd3 + 'd1)); rst_n = 'b0;
  #(100);

  if(out_valid !== 1'b0 || out_data !== 8'd0) begin : RESET_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("           Output must be 0 after reset           ");
    $display("--------------------------------------------------");
      #(CYCLE * 5);
    $finish;
  end

  #(CYCLE * 0.25); rst_n = 'b1;
  #(CYCLE); release clk;
  repeat(3) @(negedge clk);
endtask

task input_task;
  // repeat($random(SEED) % 'd3 + 'd1) @(negedge clk);
    @(negedge clk);
  // Generate random inputs
  test_pic_no = $random(SEED) % 'd16;
  test_mode = $random(SEED) % 'd2;
  test_ratio_mode = $random(SEED) % 'd4;
  // Send inputs
  in_valid = 1'b1;
  in_pic_no = test_pic_no;
  in_mode = test_mode;
  in_ratio_mode = in_mode ? test_ratio_mode : 'dx;
    @(negedge clk);
  // Reset inputs
  in_valid = 1'b0;
  in_pic_no = 'dx; in_mode = 'dx; in_ratio_mode = 'dx;
    @(negedge clk);
  exe_latency = 1;
endtask

integer contrast2_de, contrast4_de, contrast6_de;
integer adder[11:0];
task ans_gen_task;
  foreach(pic[i, j, k])
    pic[i][j][k] = DRAM[test_pic_no][i][j][k];
  case(test_mode)
    1'b0: begin
      // Auto Focus
      foreach(gray_pic[i, j])
        gray_pic[i][j] = (pic[0][i][j] >> 2) + (pic[1][i][j] >> 1) + (pic[2][i][j] >> 2);
      contrast2 = 0;
      contrast4 = 0;
      contrast6 = 0;
      foreach(gray_pic[i, j]) begin
        if(i >= 15 && i <= 16 && j >= 15 && j <= 16) begin
          if(i != 16)
            contrast2 = contrast2 + diff(gray_pic[i][j], gray_pic[i + 1][j]);
          if(j != 16)
            contrast2 = contrast2 + diff(gray_pic[i][j], gray_pic[i][j + 1]);
        end
        if(i >= 14 && i <= 17 && j >= 14 && j <= 17) begin
          if(i != 17)
            contrast4 = contrast4 + diff(gray_pic[i][j], gray_pic[i + 1][j]);
          if(j != 17)
            contrast4 = contrast4 + diff(gray_pic[i][j], gray_pic[i][j + 1]);
        end
        if(i >= 13 && i <= 18 && j >= 13 && j <= 18) begin
          if(i != 18) begin
            contrast6 = contrast6 + diff(gray_pic[i][j], gray_pic[i + 1][j]);
          end
          if(j != 18) begin
            contrast6 = contrast6 + diff(gray_pic[i][j], gray_pic[i][j + 1]);
          end
        end
      end
      contrast2_de = contrast2;
      contrast4_de = contrast4;
      contrast6_de = contrast6;
      contrast2 = contrast2 / 4;
      contrast4 = contrast4 / 16;
      contrast6 = contrast6 / 36;
      if(contrast2 >= contrast4 && contrast2 >= contrast6)
        golden_out = 8'h00;
      else if(contrast4 >= contrast2 && contrast4 >= contrast6)
        golden_out = 8'h01;
      else
        golden_out = 8'h02;
    end
    1'b1: begin
      // Auto Exposure
      case(test_ratio_mode)
        2'b00: foreach(pic[i, j, k]) pic[i][j][k] = pic[i][j][k] >> 2;
        2'b01: foreach(pic[i, j, k]) pic[i][j][k] = pic[i][j][k] >> 1;
        2'b10: foreach(pic[i, j, k]) pic[i][j][k] = pic[i][j][k];
        2'b11: foreach(pic[i, j, k]) pic[i][j][k] = pic[i][j][k][7] ? 8'hff : pic[i][j][k] << 1;
      endcase
      foreach(pic[i, j, k])
        DRAM[test_pic_no][i][j][k] = pic[i][j][k];
      expos_sum = 0;
      foreach(gray_pic[i, j]) begin
        gray_pic[i][j] = (pic[0][i][j] >> 2) + (pic[1][i][j] >> 1) + (pic[2][i][j] >> 2);
        expos_sum = expos_sum + gray_pic[i][j];
      end
      golden_out = expos_sum / 1024;
    end
  endcase
  if(`DEBUG_MODE) begin
    f_debug = $fopen("debug.txt", "w");
    $fdisplay(f_debug, "Pattern No. %4d", pat_count);
    if(test_mode) begin
      $fdisplay(f_debug, "Mode: Auto Exposure with Ratio Mode %2d", test_ratio_mode);
      $fdisplay(f_debug, "sum: %7d", expos_sum);
    end else
      $fdisplay(f_debug, "Mode: Auto Focus");
    $fdisplay(f_debug, "Picture No.: %2d", test_pic_no);
    $fdisplay(f_debug, "(R)");
    print_array(f_debug, pic[0], ~test_mode);
    $fdisplay(f_debug, "(G)");
    print_array(f_debug, pic[1], ~test_mode);
    $fdisplay(f_debug, "(B)");
    print_array(f_debug, pic[2], ~test_mode);
    $fdisplay(f_debug, "Gray Picture");
    print_array(f_debug, gray_pic, ~test_mode);
    if(test_mode == 0) begin
      $fdisplay(f_debug, "Contrast 2x2 sum: %3d", contrast2_de);
      $fdisplay(f_debug, "Contrast 4x4 sum: %3d", contrast4_de);
      $fdisplay(f_debug, "Contrast 6x6 sum: %3d", contrast6_de);
      $fdisplay(f_debug, "Contrast 2x2: %3d", contrast2);
      $fdisplay(f_debug, "Contrast 4x4: %3d", contrast4);
      $fdisplay(f_debug, "Contrast 6x6: %3d", contrast6);
    end
    $fdisplay(f_debug, "Golden Output: %3d", golden_out);
    $fclose(f_debug);
  end
endtask

function integer diff;
  input reg [7:0] a, b;
  begin
    diff = (a > b) ? (a - b) : (b - a);
  end
endfunction

task print_array;
  input integer file;
  input reg [7:0] array[0:31][0:31];
  input reg part;
  integer p, q;
  integer idx_s, idx_e;
  begin
    idx_s = part ? 13 : 0;
    idx_e = part ? 18 : 31;
    $fwrite(file, "    ");
    for(p = idx_s; p <= idx_e; p = p + 1)
      $fwrite(file, "%3d ", p);
    $fwrite(file, "\n----");
    for(p = idx_s; p <= idx_e; p = p + 1)
      $fwrite(file, "----");
    $fwrite(file, "\n");
    for(p = idx_s; p <= idx_e; p = p + 1) begin
      $fwrite(file, "%2d| ", p);
      for(q = idx_s; q <= idx_e; q = q + 1) begin
        $fwrite(file, "%3d ", array[p][q]);
      end
      $fwrite(file, "\n");
    end
    $fwrite(file, "\n");
  end
endtask

task wait_task;
  while(out_valid !== 1'b1) begin
    exe_latency = exe_latency + 1;
    if(exe_latency == 20000) begin : TIMEOUT_CHECK
      fail_task;
      $display("--------------------------------------------------");
      $display("                      FAIL!!                      ");
      $display("       Execution timeout (over 20000 cycles)       ");
      $display("--------------------------------------------------");
      repeat(5) @(negedge clk);
      $finish;
    end
      @(negedge clk);
  end
endtask

task check_task;
  rec_out = out_data;
  check = 0;
  if(test_mode === 1) begin
    check = (rec_out !== golden_out && rec_out + 1 !== golden_out && rec_out - 1 !== golden_out);
  end
  if(test_mode === 0) begin
    check = (rec_out !== golden_out);
  end
    @(negedge clk);
  if(out_valid !== 1'b0) begin
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("        out_valid must be low after output        ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
  if(check) begin
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("         Output does not match with golden        ");
    $display("==================================================\n");
    $display("  Pattern No. %4d", pat_count);
    $display("  Mode: %s", test_mode ? "Auto Exposure" : "Auto Focus");
    $display("\n  Golden Output:   %3d", golden_out);
    $display("  Received Output: %3d", rec_out);
    $display("\n--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
  $display("\033[38;5;123mPATTERN NO.%4d PASS!!\033[0;32m EXECUTION CYCLE :%4d\033[m", pat_count, exe_latency);
  total_latency = total_latency + exe_latency;
endtask

//================================================================
// ASCII Art
//================================================================
task YOU_PASS_task;
  $display("[38;2;0;0;0m                                          [38;2;0;1;0m [38;2;5;2;5m [38;2;17;6;13m'[38;2;32;13;25m,[38;2;55;19;40ml[38;2;73;22;52mi[38;2;92;22;64m+[38;2;98;20;66m_[38;2;99;19;65m_[38;2;102;19;66m_[38;2;105;19;67m_[38;2;103;20;67m_[38;2;101;19;66m_[38;2;101;17;65m_[38;2;102;16;64m_[38;2;102;17;65m_[38;2;101;18;65m_[38;2;99;18;64m_______________[38;2;101;18;65m_[38;2;102;18;65m_[38;2;103;19;67m__[38;2;102;20;67m_[38;2;104;21;65m_[38;2;94;23;60m+[38;2;65;17;42ml[38;2;30;10;19m\"[38;2;5;2;3m [38;2;0;0;0m                                                                                          [38;2;0;0;0m");
  $display("[38;2;0;0;0m                                        [38;2;10;4;8m.[38;2;36;11;27m,[38;2;64;17;44ml[38;2;89;18;58m+[38;2;103;20;69m-[38;2;108;22;73m-[38;2;113;20;75m?[38;2;116;18;75m?[38;2;115;18;73m-[38;2;114;17;73m-[38;2;114;18;73m--[38;2;115;18;73m-[38;2;114;18;73m-[38;2;111;18;72m-[38;2;111;17;71m-[38;2;112;16;71m-[38;2;111;17;71m-[38;2;110;18;71m-[38;2;110;17;71m--------------[38;2;110;17;72m---[38;2;111;18;73m--[38;2;112;18;73m-[38;2;115;18;73m-[38;2;118;18;74m?[38;2;119;18;74m?[38;2;113;20;69m-[38;2;88;22;57m+[38;2;49;14;34mI[38;2;12;4;9m.[38;2;0;0;0m                                                                                        [38;2;0;0;0m");
  $display("[38;2;0;0;0m                                 [38;2;0;0;1m  [38;2;0;1;0m [38;2;0;0;0m  [38;2;22;8;14m^[38;2;59;17;41ml[38;2;92;21;63m+[38;2;111;20;72m-[38;2;115;19;73m?[38;2;114;18;73m-[38;2;112;18;73m-[38;2;112;18;72m-[38;2;111;17;71m-[38;2;111;17;70m-[38;2;111;18;70m---[38;2;111;17;70m-[38;2;111;18;70m--[38;2;110;17;70m----------------[38;2;110;18;69m-[38;2;109;18;70m-[38;2;109;18;71m-[38;2;109;18;72m-[38;2;110;17;71m--[38;2;111;18;72m--[38;2;110;18;73m-[38;2;112;17;74m-[38;2;113;17;73m-[38;2;113;18;73m-[38;2;116;18;73m?[38;2;119;17;73m?[38;2;115;21;75m?[38;2;94;24;64m_[38;2;55;17;37mI[38;2;16;7;11m'[38;2;0;1;0m [38;2;0;0;0m                                                                                     [38;2;0;0;0m");
  $display("[38;2;0;0;0m                                    [38;2;21;6;12m'[38;2;63;17;43ml[38;2;103;21;68m-[38;2;117;17;74m?[38;2;113;17;72m-[38;2;111;17;71m--[38;2;111;18;71m-[38;2;111;18;70m-[38;2;111;18;71m-[38;2;110;17;70m-----------------------[38;2;110;17;71m-[38;2;111;18;70m-[38;2;112;18;71m-[38;2;112;16;73m-[38;2;112;16;74m-[38;2;110;16;71m-[38;2;109;15;68m-[38;2;108;16;67m_[38;2;107;17;65m_[38;2;107;19;63m_[38;2;107;18;66m_[38;2;108;16;69m-[38;2;109;16;71m-[38;2;113;17;72m-[38;2;115;17;72m-[38;2;111;19;72m-[38;2;112;19;74m-[38;2;113;20;75m?[38;2;94;23;64m_[38;2;57;19;41ml[38;2;20;7;17m^[38;2;0;1;3m [38;2;0;0;0m                                                                                   [38;2;0;0;0m");
  $display("[38;2;0;0;0m                              [38;2;1;0;0m [38;2;0;0;0m   [38;2;14;5;8m.[38;2;56;16;35mI[38;2;101;21;64m_[38;2;116;19;73m?[38;2;115;16;73m-[38;2;112;17;71m-[38;2;111;18;70m-[38;2;110;17;70m---------------------------[38;2;111;17;67m-[38;2;110;16;68m-[38;2;110;15;69m-[38;2;108;13;66m_[38;2;105;16;62m_[38;2;104;27;59m_[38;2;109;41;59m?[38;2;119;62;63mt[38;2;125;82;62mj[38;2;132;99;64mx[38;2;137;109;66mn[38;2;136;104;67mn[38;2;126;82;62mj[38;2;115;59;59m1[38;2;109;40;61m?[38;2;107;26;63m-[38;2;107;20;66m-[38;2;108;18;68m-[38;2;110;17;72m-[38;2;111;18;74m-[38;2;112;21;71m-[38;2;101;22;68m_[38;2;66;18;48m![38;2;25;9;21m^[38;2;3;2;3m [38;2;0;0;0m [38;2;0;0;1m [38;2;2;0;1m [38;2;1;0;0m [38;2;0;0;0m                                                                             [38;2;0;0;0m");
  $display("[38;2;0;0;0m                             [38;2;1;0;0m [38;2;2;0;0m [38;2;0;1;0m [38;2;4;1;1m [38;2;42;12;27m,[38;2;92;23;60m+[38;2;116;19;71m-[38;2;113;17;70m--[38;2;113;17;71m-[38;2;110;17;70m------------------------[38;2;111;18;71m--[38;2;112;17;72m-[38;2;110;16;72m-[38;2;106;13;67m_[38;2;107;16;61m_[38;2;111;34;62m?[38;2;123;63;69mf[38;2;145;101;79mu[38;2;161;135;83mX[38;2;174;160;86mJ[38;2;183;170;95mL[38;2;167;155;81mU[38;2;156;146;71mX[38;2;155;146;72mX[38;2;169;161;84mJ[38;2;175;164;84mJ[38;2;158;148;70mX[38;2;151;142;72mz[38;2;141;129;67mv[38;2;138;119;68mu[38;2;130;99;63mx[38;2;118;74;58mf[38;2;109;52;57m?[38;2;106;32;60m-[38;2;107;21;64m-[38;2;107;19;70m-[38;2;111;21;73m-[38;2;105;23;71m-[38;2;82;20;58m~[38;2;43;15;31m;[38;2;13;6;9m.[38;2;0;1;0m [38;2;0;0;0m                                                                              [38;2;0;0;0m");
  $display("[38;2;0;0;0m                             [38;2;1;0;1m [38;2;0;1;0m [38;2;11;4;7m.[38;2;66;18;43m![38;2;107;21;69m-[38;2;112;17;71m-[38;2;111;17;70m-[38;2;110;17;69m-[38;2;110;17;70m----------------------[38;2;111;17;70m-[38;2;109;18;70m-[38;2;108;18;71m-[38;2;112;17;72m-[38;2;112;16;74m-[38;2;109;14;73m-[38;2;105;19;65m_[38;2;112;39;64m?[38;2;138;81;77mx[38;2;171;137;92mU[38;2;199;185;107mO[38;2;213;208;117mq[38;2;218;216;119mp[38;2;217;216;117mp[38;2;213;212;117mq[38;2;210;208;117mw[38;2;205;202;109mm[38;2;162;155;72mY[38;2;136;126;57mu[38;2;184;176;99mQ[38;2;216;210;120mq[38;2;196;191;99mO[38;2;163;157;76mY[38;2;138;130;60mu[38;2;176;172;87mC[38;2;175;172;82mC[38;2;161;156;75mY[38;2;153;143;69mz[38;2;147;127;69mv[38;2;138;109;68mn[38;2;125;80;63mj[38;2;109;45;60m?[38;2;103;22;59m_[38;2;111;19;76m-[38;2;112;22;75m?[38;2;99;23;63m_[38;2;67;19;42m![38;2;28;9;17m^[38;2;2;1;0m [38;2;0;1;0m [38;2;0;1;1m [38;2;0;0;0m                                                                          [38;2;0;0;0m");
  $display("[38;2;0;0;0m                              [38;2;18;6;12m'[38;2;84;21;55m~[38;2;112;20;72m-[38;2;111;17;70m-[38;2;110;17;70m---------------------[38;2;111;17;70m-[38;2;113;16;70m-[38;2;110;17;70m-[38;2;106;17;68m_[38;2;106;15;68m_[38;2;109;15;70m-[38;2;109;17;69m-[38;2;102;17;64m_[38;2;102;26;60m_[38;2;119;67;64mf[38;2;159;133;87mX[38;2;200;188;115mZ[38;2;216;211;121mq[38;2;215;216;119mp[38;2;213;213;114mq[38;2;213;210;111mw[38;2;213;211;111mw[38;2;214;211;115mq[38;2;189;185;99m0[38;2;200;196;109mZ[38;2;217;213;120mp[38;2;177;170;87mC[38;2;134;124;55mn[38;2;200;193;111mZ[38;2;214;211;113mq[38;2;216;212;111mq[38;2;207;202;114mw[38;2;160;152;78mY[38;2;209;204;113mw[38;2;216;212;115mq[38;2;206;201;113mm[38;2;175;170;88mC[38;2;167;161;85mU[38;2;150;145;68mz[38;2;145;140;62mc[38;2;151;135;75mz[38;2;125;91;60mr[38;2;100;45;58m-[38;2;99;23;61m_[38;2;109;17;73m-[38;2;116;19;77m?[38;2;107;22;67m-[38;2;70;19;46m![38;2;23;7;15m^[38;2;0;0;0m                               [38;2;3;4;2m [38;2;19;21;19m\"[38;2;15;17;15m^[38;2;0;0;0m                                         [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;1;0;0m [38;2;1;0;1m [38;2;0;1;0m [38;2;0;0;0m [38;2;22;7;14m^[38;2;88;22;56m+[38;2;114;16;72m-[38;2;110;17;69m-[38;2;109;18;68m-[38;2;110;17;70m--------------[38;2;108;18;70m-[38;2;109;18;70m-[38;2;111;17;70m--[38;2;110;17;70m--[38;2;111;17;70m-[38;2;109;17;71m-[38;2;106;15;68m_[38;2;102;13;63m+[38;2;103;14;67m_[38;2;107;16;70m-[38;2;105;16;72m-[38;2;107;35;65m?[38;2;129;84;65mr[38;2;176;157;96mC[38;2;213;205;116mw[38;2;221;219;117mp[38;2;202;201;105mZ[38;2;191;191;98mO[38;2;211;212;116mq[38;2;210;211;111mw[38;2;211;211;110mw[38;2;208;207;113mw[38;2;189;186;100m0[38;2;193;190;107mO[38;2;213;210;119mq[38;2;215;211;123mp[38;2;163;158;76mY[38;2;176;171;88mC[38;2;216;212;117mq[38;2;215;211;113mq[38;2;212;208;115mw[38;2;188;183;94mQ[38;2;197;192;103mO[38;2;215;211;117mq[38;2;213;210;114mq[38;2;214;212;115mq[38;2;196;194;109mZ[38;2;215;212;148md[38;2;190;190;113mO[38;2;138;133;57mu[38;2;161;155;76mY[38;2;169;161;78mU[38;2;152;135;76mz[38;2;129;98;65mx[38;2;105;51;59m?[38;2;99;21;64m_[38;2;109;19;73m-[38;2;114;22;77m?[38;2;102;25;69m-[38;2;39;14;24m,[38;2;1;0;0m  [38;2;0;0;0m [38;2;1;0;0m [38;2;0;0;0m                         [38;2;18;21;18m\"[38;2;158;167;157mO[38;2;199;203;195mk[38;2;208;212;203ma[38;2;109;112;106mu[38;2;0;0;0m  [38;2;0;0;2m [38;2;0;0;0m                                     [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;1;0;1m [38;2;0;0;0m [38;2;11;3;8m.[38;2;83;22;54m~[38;2;117;18;71m-[38;2;115;16;71m-[38;2;110;17;69m-[38;2;112;16;70m-[38;2;110;17;70m--------------[38;2;108;18;70m-[38;2;109;18;70m-[38;2;111;17;70m---[38;2;108;17;70m-[38;2;101;14;65m_[38;2;94;11;60m+[38;2;98;13;63m+[38;2;105;16;67m_[38;2;102;21;66m_[38;2;102;39;60m-[38;2;128;89;70mr[38;2;173;158;92mJ[38;2;209;209;115mw[38;2;221;218;118mp[38;2;213;209;112mw[38;2;195;193;103mO[38;2;188;186;99m0[38;2;209;208;115mw[38;2;214;213;119mq[38;2;210;209;115mw[38;2;198;196;105mZ[38;2;187;184;107m0[38;2;223;219;151mk[38;2;231;228;151mh[38;2;212;208;119mq[38;2;190;185;101m0[38;2;190;185;103m0[38;2;226;222;132mb[38;2;213;213;114mq[38;2;202;199;111mm[38;2;170;166;86mJ[38;2;188;185;100m0[38;2;225;221;128md[38;2;213;209;119mq[38;2;216;213;123mp[38;2;216;215;118mp[38;2;205;205;115mw[38;2;202;200;134mw[38;2;234;235;163ma[38;2;182;182;99mQ[38;2;180;178;95mQ[38;2;214;212;118mq[38;2;197;193;107mZ[38;2;171;168;82mJ[38;2;151;139;70mz[38;2;127;90;65mr[38;2;102;36;54m-[38;2;110;22;69m-[38;2;120;19;76m?[38;2;99;29;60m_[38;2;27;11;15m^[38;2;0;0;0m  [38;2;2;0;0m [38;2;0;0;0m                         [38;2;24;25;23m,[38;2;165;168;157mO[38;2;174;175;158mZ[38;2;206;210;196mh[38;2;149;153;147mL[38;2;0;0;0m  [38;2;0;0;2m [38;2;0;0;0m                                     [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;1;1;0m [38;2;1;0;0m [38;2;41;14;32m;[38;2;95;15;60m+[38;2;97;11;61m+[38;2;102;14;63m+[38;2;110;17;68m-[38;2;112;17;70m-[38;2;111;17;70m-[38;2;109;17;70m-[38;2;108;18;70m-[38;2;110;17;70m-----------[38;2;109;17;70m-[38;2;110;17;70m-[38;2;112;17;70m-[38;2;113;17;70m-[38;2;105;17;67m_[38;2;93;10;59m~[38;2;93;10;58m~[38;2;103;14;66m_[38;2;107;18;66m_[38;2;104;33;61m-[38;2;122;81;65mj[38;2;157;140;79mX[38;2;200;194;108mZ[38;2;214;212;116mq[38;2;200;197;109mZ[38;2;175;170;86mC[38;2;168;164;79mU[38;2;197;193;106mZ[38;2;227;225;140mk[38;2;227;226;145mk[38;2;200;200;117mm[38;2;184;186;105m0[38;2;205;206;131mq[38;2;244;243;180m#[38;2;252;250;187mW[38;2;212;211;128mp[38;2;188;186;97m0[38;2;201;198;112mm[38;2;224;222;135mb[38;2;205;203;115mw[38;2;192;191;104mO[38;2;189;187;106mO[38;2;182;180;97mQ[38;2;219;218;127md[38;2;217;216;121mp[38;2;207;205;115mw[38;2;191;189;104mO[38;2;221;221;128md[38;2;208;209;117mw[38;2;193;193;124mm[38;2;234;235;165mo[38;2;193;192;107mO[38;2;196;195;109mZ[38;2;214;213;119mq[38;2;213;212;114mq[38;2;213;210;117mq[38;2;194;191;102mO[38;2;163;156;79mY[38;2;133;109;65mn[38;2;106;35;56m-[38;2;112;19;73m-[38;2;111;22;73m-[38;2;73;19;47mi[38;2;4;1;3m [38;2;0;0;0m [38;2;0;1;0m [38;2;0;0;0m                         [38;2;21;21;20m\"[38;2;153;156;145mQ[38;2;169;173;151mO[38;2;200;204;186mb[38;2;140;142;136mJ[38;2;0;0;0m                                        [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;1;0;0m [38;2;0;0;0m [38;2;8;3;4m.[38;2;65;15;41ml[38;2;83;8;50mi[38;2;80;7;48m![38;2;83;7;50mi[38;2;91;12;55m~[38;2;105;18;68m_[38;2;109;17;70m-[38;2;110;17;70m---------------[38;2;109;19;71m-[38;2;105;15;67m_[38;2;96;10;59m+[38;2;102;12;63m+[38;2;108;19;70m-[38;2;105;20;66m_[38;2;118;57;59mt[38;2;146;122;73mv[38;2;159;153;81mY[38;2;187;180;99mQ[38;2;183;175;96mQ[38;2;162;156;78mY[38;2;148;143;68mz[38;2;165;163;85mU[38;2;210;208;129mq[38;2;228;226;149mk[38;2;214;211;134mp[38;2;192;192;109mO[38;2;204;205;125mw[38;2;233;234;165ma[38;2;250;251;189mW[38;2;234;235;169mo[38;2;196;196;118mm[38;2;185;185;97mQ[38;2;197;196;108mZ[38;2;201;198;112mm[38;2;197;195;108mZ[38;2;198;196;110mZ[38;2;195;193;107mZ[38;2;188;186;100m0[38;2;208;207;113mw[38;2;212;212;114mq[38;2;207;207;112mw[38;2;206;205;114mw[38;2;179;177;92mL[38;2;212;211;119mq[38;2;209;208;114mw[38;2;190;188;112mO[38;2;213;213;134mp[38;2;178;176;91mL[38;2;214;213;120mq[38;2;213;214;115mq[38;2;210;209;110mw[38;2;212;210;111mw[38;2;216;214;115mq[38;2;205;202;110mm[38;2;164;158;82mU[38;2;105;70;54m1[38;2;102;20;59m_[38;2;115;20;71m-[38;2;84;24;56m~[38;2;7;2;5m [38;2;0;0;0m [38;2;0;1;0m [38;2;0;0;0m                         [38;2;19;19;18m^[38;2;154;156;145mQ[38;2;172;175;156mZ[38;2;207;208;196mh[38;2;139;139;138mJ[38;2;0;0;0m                                        [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;0;1;0m [38;2;21;9;17m^[38;2;75;13;47m![38;2;79;9;50mi[38;2;79;8;48m![38;2;82;8;49mi[38;2;83;7;48mi[38;2;92;11;56m~[38;2;106;19;69m-[38;2;109;18;70m-[38;2;110;17;72m-[38;2;110;17;70m------------[38;2;109;17;70m-[38;2;105;16;68m_[38;2;98;9;61m+[38;2;104;16;67m_[38;2;109;21;69m-[38;2;107;18;68m-[38;2;107;45;61m?[38;2;156;132;78mz[38;2;155;149;67mz[38;2;155;144;73mX[38;2;155;143;69mz[38;2;146;137;68mc[38;2;154;147;75mX[38;2;188;184;101m0[38;2;202;201;118mm[38;2;201;199;116mm[38;2;198;196;111mZ[38;2;202;201;112mm[38;2;216;217;124mp[38;2;234;234;151ma[38;2;221;220;143mb[38;2;195;195;118mZ[38;2;180;180;98mQ[38;2;184;185;97mQ[38;2;193;194;104mO[38;2;196;195;101mO[38;2;205;204;112mm[38;2;200;198;112mm[38;2;187;184;100m0[38;2;194;192;103mO[38;2;210;210;116mw[38;2;211;211;111mw[38;2;214;214;113mq[38;2;193;190;97mO[38;2;190;186;99m0[38;2;185;181;95mQ[38;2;215;212;118mq[38;2;201;197;105mZ[38;2;188;184;98m0[38;2;189;186;97m0[38;2;206;203;112mm[38;2;214;212;117mq[38;2;212;210;111mw[38;2;210;209;111mw[38;2;210;210;111mw[38;2;211;211;112mw[38;2;213;213;114mq[38;2;213;212;117mq[38;2;161;153;89mU[38;2;106;50;58m?[38;2;109;21;68m-[38;2;84;22;54m~[38;2;5;1;4m [38;2;0;1;0m [38;2;1;1;0m [38;2;0;0;0m                         [38;2;15;16;14m^[38;2;108;112;105mu[38;2;118;120;114mc[38;2;191;191;189md[38;2;136;136;136mU[38;2;0;0;0m                                        [38;2;0;0;0m");
  $display("[38;2;0;0;0m                           [38;2;30;12;24m\"[38;2;80;13;49mi[38;2;77;10;50m![38;2;78;10;49m![38;2;80;9;49mi[38;2;81;9;49mi[38;2;83;6;49mi[38;2;96;12;60m+[38;2;109;18;70m-[38;2;113;15;72m-[38;2;110;17;70m------------[38;2;109;18;70m-[38;2;102;13;65m_[38;2;104;15;66m_[38;2;111;19;70m-[38;2;108;20;70m-[38;2;100;26;57m_[38;2;134;103;71mn[38;2;156;146;74mX[38;2;151;142;67mz[38;2;155;142;71mz[38;2;149;137;67mc[38;2;171;163;91mJ[38;2;193;188;108mO[38;2;199;196;107mZ[38;2;201;200;107mZ[38;2;209;209;112mw[38;2;214;214;115mq[38;2;211;211;113mw[38;2;200;198;108mZ[38;2;181;177;95mQ[38;2;175;172;90mC[38;2;188;185;99m0[38;2;200;197;109mZ[38;2;207;205;114mw[38;2;211;210;115mw[38;2;212;212;115mq[38;2;206;206;112mw[38;2;203;202;111mm[38;2;208;207;117mw[38;2;212;212;117mq[38;2;211;211;115mq[38;2;212;213;114mq[38;2;202;200;108mm[38;2;168;162;85mJ[38;2;181;175;99mQ[38;2;208;204;112mw[38;2;214;211;114mq[38;2;196;193;101mO[38;2;207;203;112mw[38;2;210;207;110mw[38;2;215;212;113mq[38;2;206;202;110mm[38;2;204;201;108mm[38;2;212;211;112mw[38;2;210;210;112mww[38;2;211;211;113mw[38;2;212;214;112mq[38;2;204;208;113mw[38;2;129;92;69mx[38;2;105;22;67m-[38;2;74;19;50mi[38;2;2;0;2m [38;2;2;1;0m [38;2;1;1;0m [38;2;0;0;0m                         [38;2;12;13;13m'[38;2;81;85;83mf[38;2;86;88;88mj[38;2;164;164;167mZ[38;2;135;135;136mU[38;2;0;0;0m                                        [38;2;0;0;0m");
  $display("[38;2;0;0;0m                           [38;2;34;13;29m,[38;2;78;12;51mi[38;2;81;9;50mi[38;2;79;9;49m!![38;2;80;9;49mi[38;2;81;8;49mi[38;2;86;7;53mi[38;2;103;15;65m_[38;2;112;16;71m-[38;2;111;17;72m-[38;2;111;18;72m---[38;2;111;18;71m--[38;2;110;17;70m-----[38;2;110;18;69m-[38;2;110;17;70m-[38;2;109;17;71m-[38;2;110;18;73m-[38;2;113;18;69m-[38;2;108;17;68m-[38;2;113;56;67mt[38;2;154;137;77mz[38;2;154;146;67mz[38;2;175;167;84mC[38;2;200;193;104mZ[38;2;200;195;105mZ[38;2;209;205;114mw[38;2;213;210;116mq[38;2;216;214;118mq[38;2;218;217;118mp[38;2;209;207;111mw[38;2;204;201;110mm[38;2;203;200;106mZ[38;2;191;187;96m0[38;2;201;197;105mZ[38;2;213;208;120mq[38;2;184;178;100mQ[38;2;167;161;85mU[38;2;218;215;118mp[38;2;217;213;123mp[38;2;169;162;91mJ[38;2;185;181;97mQ[38;2;197;193;109mZ[38;2;185;181;96mQ[38;2;216;214;120mp[38;2;208;206;114mw[38;2;185;181;96mQ[38;2;148;142;71mz[38;2;153;143;95mY[38;2;152;141;96mY[38;2;209;203;123mw[38;2;193;188;106mO[38;2;138;130;66mv[38;2;172;167;89mC[38;2;207;203;112mw[38;2;217;214;120mp[38;2;185;180;97mQ[38;2;199;194;109mZ[38;2;211;208;114mw[38;2;212;212;116mq[38;2;212;212;112mww[38;2;214;214;116mq[38;2;212;213;124mp[38;2;132;90;70mx[38;2;109;21;68m-[38;2;64;17;41ml[38;2;1;0;0m [38;2;1;1;0m [38;2;1;0;0m [38;2;0;0;0m                         [38;2;13;15;14m^[38;2;83;87;86mf[38;2;88;89;89mj[38;2;177;174;176mw[38;2;138;136;137mU[38;2;0;0;0m                  [38;2;1;1;0m [38;2;0;0;0m     [38;2;0;1;0m [38;2;0;0;0m               [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;1;1;1m [38;2;44;14;35m;[38;2;80;10;51mi[38;2;81;9;50mi[38;2;80;9;49miii[38;2;81;8;49mi[38;2;84;7;51mi[38;2;92;8;57m~[38;2;103;15;67m_[38;2;107;13;66m___[38;2;108;14;67m_[38;2;112;18;71m-[38;2;112;19;72m-[38;2;111;18;71m--[38;2;110;17;70m---[38;2;110;18;69m-[38;2;110;17;70m-[38;2;110;17;72m-[38;2;111;18;73m-[38;2;112;18;72m-[38;2;100;23;58m_[38;2;140;104;71mn[38;2;175;167;86mC[38;2;198;195;102mZ[38;2;214;212;111mq[38;2;217;214;116mq[38;2;214;211;118mq[38;2;191;187;97m0[38;2;192;189;99mO[38;2;209;206;117mw[38;2;186;179;112m0[38;2;149;138;93mX[38;2;191;185;109mO[38;2;213;210;116mq[38;2;200;196;107mZ[38;2;179;173;97mL[38;2;156;145;99mU[38;2;137;124;86mc[38;2;185;178;106m0[38;2;198;193;111mZ[38;2;157;148;90mY[38;2;130;120;68mu[38;2;169;161;98mC[38;2;143;136;71mc[38;2;194;189;108mO[38;2;184;178;98mQ[38;2;157;150;81mY[38;2;133;122;76mv[38;2;135;121;95mc[38;2;169;153;140mQ[38;2;176;160;141m0[38;2;164;154;103mJ[38;2;166;153;115mC[38;2;187;172;150mZ[38;2;146;136;81mz[38;2;170;164;85mJ[38;2;183;176;104mQ[38;2;141;135;62mv[38;2;192;187;106mO[38;2;166;162;74mU[38;2;189;185;97m0[38;2;209;205;111mw[38;2;208;204;111mw[38;2;196;192;101mO[38;2;188;172;111m0[38;2;103;37;54m-[38;2;112;24;71m?[38;2;50;15;31mI[38;2;0;0;0m                            [38;2;19;19;19m\"[38;2;86;87;87mf[38;2;89;89;89mj[38;2;182;182;182mq[38;2;140;139;139mJ[38;2;0;0;0m                   [38;2;38;39;37ml[38;2;114;119;114mc[38;2;72;77;74m1[38;2;11;14;12m'[38;2;0;2;1m [38;2;0;0;0m                [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;4;3;3m [38;2;52;16;39mI[38;2;81;9;51mi[38;2;80;9;50mi[38;2;80;9;49miii[38;2;80;9;48m![38;2;76;6;47m![38;2;83;20;57m~[38;2;132;79;107mu[38;2;167;119;139mJ[38;2;173;130;148mL[38;2;173;126;145mL[38;2;143;84;110mv[38;2;104;25;69m-[38;2;111;20;73m-[38;2;113;19;73m-[38;2;112;19;71m-[38;2;111;18;71m-[38;2;110;17;70m----[38;2;113;18;72m-[38;2;115;19;72m-[38;2;109;18;72m-[38;2;116;57;69mt[38;2;199;184;108mO[38;2;213;212;116mq[38;2;216;214;115mq[38;2;207;204;107mm[38;2;181;176;97mQ[38;2;146;138;78mz[38;2;137;127;69mv[38;2;169;157;103mC[38;2;153;139;98mY[38;2;143;127;103mX[38;2;142;129;92mz[38;2;163;155;90mU[38;2;150;143;81mX[38;2;143;133;96mX[38;2;148;132;116mY[38;2;142;126;105mX[38;2;154;142;95mY[38;2;163;153;99mJ[38;2;152;139;108mU[38;2;135;121;93mc[38;2;137;125;85mc[38;2;136;123;89mc[38;2;138;127;82mc[38;2;152;142;86mX[38;2;139;126;85mc[38;2;150;135;110mY[38;2;166;149;138mQ[38;2;180;162;158mZ[38;2;207;191;186mb[38;2;192;177;169mq[38;2;141;127;112mX[38;2;205;189;181md[38;2;220;205;195ma[38;2;142;133;98mX[38;2;147;139;84mz[38;2;168;155;119mL[38;2;146;133;85mz[38;2;160;151;79mY[38;2;138;128;61mu[38;2;154;147;74mX[38;2;168;162;84mJ[38;2;182;176;99mQ[38;2;161;154;83mY[38;2;120;82;62mj[38;2;101;19;64m_[38;2;110;27;71m?[38;2;36;12;21m,[38;2;0;0;0m [38;2;0;1;0m [38;2;0;0;0m                       [38;2;0;0;1m [38;2;2;0;0m [38;2;36;33;32mI[38;2;65;66;63m-[38;2;88;86;89mj[38;2;91;89;93mj[38;2;186;185;186mp[38;2;193;192;191mb[38;2;127;126;124mX[38;2;48;48;46mi[38;2;0;0;0m  [38;2;18;18;19m^[38;2;41;41;44m![38;2;46;46;49mi[38;2;49;50;53mi[38;2;51;52;56m~[38;2;53;54;59m+[38;2;58;58;65m_[38;2;62;64;71m-[38;2;67;69;75m?[38;2;70;72;78m?[38;2;72;75;81m1[38;2;75;78;84mt[38;2;78;81;87mt[38;2;87;90;96mj[38;2;100;102;108mn[38;2;115;118;123mc[38;2;165;170;175mm[38;2;174;180;183mq[38;2;136;142;148mC[38;2;122;129;135mY[38;2;39;45;42m![38;2;0;0;0m    [38;2;0;0;1m    [38;2;0;0;0m       [38;2;0;0;0m");
  $display("[38;2;33;34;32mI[38;2;36;36;35mI[38;2;37;37;36mI[38;2;38;39;37ml[38;2;41;41;39ml[38;2;42;42;41mll[38;2;43;43;41m![38;2;41;41;39ml[38;2;39;38;35ml[38;2;36;36;33mI[38;2;41;41;38ml[38;2;45;45;42m![38;2;49;49;46mi[38;2;51;50;48mi[38;2;52;53;52m~[38;2;53;54;53m~[38;2;55;56;55m+[38;2;57;57;56m+[38;2;59;59;58m+[38;2;59;59;59m+[38;2;61;62;61m_[38;2;61;63;60m_[38;2;60;63;60m_[38;2;56;59;56m+[38;2;7;9;7m.[38;2;5;3;4m [38;2;60;17;42ml[38;2;85;7;51mi[38;2;78;9;49m![38;2;80;9;49mi[38;2;80;9;50mi[38;2;80;9;49mi[38;2;76;7;45m![38;2;90;36;61m_[38;2;193;160;167mm[38;2;228;211;205mo[38;2;227;215;205m*[38;2;226;216;204m*[38;2;229;216;206m*[38;2;231;211;206m*[38;2;149;103;122mX[38;2;103;20;64m_[38;2;118;19;75m?[38;2;114;20;74m?[38;2;111;18;71m-[38;2;110;17;70m----[38;2;113;18;71m-[38;2;116;18;74m?[38;2;102;20;60m_[38;2;169;130;100mU[38;2;217;210;123mp[38;2;201;198;106mZ[38;2;186;180;100mQ[38;2;148;137;87mX[38;2;144;130;103mX[38;2;126;113;90mu[38;2;127;116;92mv[38;2;141;129;115mY[38;2;145;132;128mU[38;2;132;120;110mz[38;2;143;134;120mY[38;2;145;137;128mU[38;2;147;139;135mJ[38;2;147;136;134mJ[38;2;132;117;114mz[38;2;136;120;104mz[38;2;161;146;126mC[38;2;171;154;146m0[38;2;139;122;118mX[38;2;144;127;115mY[38;2;176;160;147mO[38;2;187;170;166mw[38;2;138;122;107mz[38;2;153;136;124mU[38;2;187;168;163mmm[38;2;160;142;138mC[38;2;156;143;142mL[38;2;175;168;172mm[38;2;183;179;186mq[38;2;192;191;202mb[38;2;204;202;211mh[38;2;199;198;206mk[38;2;164;162;166mO[38;2;147;139;136mJ[38;2;172;157;152mO[38;2;149;135;108mY[38;2;129;117;68mn[38;2;143;133;67mv[38;2;155;146;72mX[38;2;154;145;72mz[38;2;143;133;67mv[38;2;154;141;85mX[38;2;93;47;45m_[38;2;105;23;71m-[38;2;105;29;66m-[38;2;25;9;14m^[38;2;0;0;0m           [38;2;2;2;4m [38;2;28;27;30m;[38;2;40;39;42ml[38;2;62;61;65m_[38;2;94;94;97mr[38;2;97;99;102mx[38;2;88;90;94mj[38;2;76;75;81m1[38;2;77;77;80mt[38;2;57;57;58m+[38;2;2;3;3m [38;2;0;0;0m    [38;2;42;37;39ml[38;2;96;91;94mr[38;2;85;85;86mf[38;2;88;86;89mj[38;2;92;90;96mr[38;2;194;192;193mb[38;2;195;196;189mb[38;2;175;177;165mm[38;2;191;191;180mp[38;2;85;81;76mt[38;2;59;52;53m~[38;2;116;110;114mv[38;2;163;162;169mO[38;2;155;157;167m0[38;2;153;155;167m0[38;2;152;155;168m0[38;2;152;154;169m0[38;2;151;154;169m0[38;2;148;153;166mQ[38;2;147;152;164mQ[38;2;145;150;162mQ[38;2;146;148;160mQ[38;2;145;146;157mL[38;2;144;145;157mL[38;2;142;142;154mC[38;2;139;139;152mC[38;2;133;133;146mU[38;2;124;124;137mY[38;2;123;123;135mX[38;2;130;131;149mU[38;2;154;160;172mO[38;2;56;62;58m+[38;2;0;0;0m [38;2;0;1;1m [38;2;1;2;2m [38;2;2;3;3m  [38;2;3;3;3m [38;2;5;4;4m [38;2;8;5;5m.[38;2;9;6;6m.[38;2;10;8;7m.[38;2;11;9;8m..[38;2;12;9;9m'[38;2;12;10;10m'[38;2;13;11;10m'[38;2;14;12;10m'");
  $display("[38;2;179;181;169mww[38;2;180;182;169mw[38;2;181;183;169mww[38;2;180;183;169mw[38;2;181;182;168mw[38;2;177;170;159mZ[38;2;192;182;173mq[38;2;204;192;183mb[38;2;205;192;184mb[38;2;209;196;187mk[38;2;190;180;171mq[38;2;181;176;165mw[38;2;188;188;176mp[38;2;187;191;179mp[38;2;189;191;180mp[38;2;190;193;181md[38;2;191;193;182md[38;2;192;194;182md[38;2;193;196;183md[38;2;195;197;185mb[38;2;195;198;186mb[38;2;196;201;188mb[38;2;203;207;197mh[38;2;45;50;46mi[38;2;11;4;7m.[38;2;71;17;45m![38;2;83;9;48mi[38;2;80;9;47m!![38;2;81;10;48mi[38;2;81;10;49mi[38;2;73;10;42ml[38;2;156;118;129mU[38;2;236;214;208m*[38;2;223;207;201ma[38;2;224;206;199ma[38;2;225;206;199ma[38;2;225;207;198ma[38;2;229;213;203m*[38;2;201;171;176mq[38;2;109;31;71m?[38;2;120;17;74m?[38;2;116;19;73m?[38;2;112;18;71m-[38;2;108;18;70m-[38;2;109;17;70m-[38;2;110;17;70m--[38;2;112;19;72m-[38;2;113;19;73m-[38;2;108;35;63m-[38;2;175;149;118mL[38;2;155;143;95mY[38;2;149;139;91mX[38;2;132;120;88mv[38;2;149;137;130mJ[38;2;167;158;160mO[38;2;151;151;153mQ[38;2;174;178;183mw[38;2;199;202;211mh[38;2;205;207;217ma[38;2;207;209;221mo[38;2;216;219;229m#[38;2;215;220;230m#[38;2;210;215;226m*[38;2;187;187;193md[38;2;147;138;137mJ[38;2;154;136;134mJ[38;2;180;160;158mZ[38;2;181;163;159mZ[38;2;148;129;126mU[38;2;147;129;124mU[38;2;203;185;178md[38;2;220;201;196mh[38;2;195;177;170mq[38;2;204;185;180md[38;2;195;176;170mq[38;2;146;134;131mU[38;2;174;170;173mm[38;2;226;229;234mW[38;2;232;234;238m&[38;2;184;179;185mq[38;2;243;241;247mB[38;2;245;245;249mB[38;2;244;246;252m@[38;2;229;227;237mW[38;2;107;96;109mn[38;2;116;101;100mn[38;2;163;147;138mL[38;2;173;158;134mQ[38;2;147;136;74mz[38;2;157;145;70mX[38;2;153;137;77mz[38;2;112;83;54mf[38;2;138;110;77mu[38;2;121;78;67mj[38;2;104;27;66m-[38;2;101;29;63m-[38;2;26;12;15m^[38;2;12;9;7m.[38;2;14;10;8m'[38;2;17;11;9m'[38;2;20;15;11m^[38;2;22;17;13m^[38;2;23;18;14m^[38;2;27;21;16m\"[38;2;30;22;18m,[38;2;30;24;20m,[38;2;32;26;21m,[38;2;36;29;26m;[38;2;77;73;76m1[38;2;139;139;150mC[38;2;139;139;153mC[38;2;139;141;153mC[38;2;139;142;154mC[38;2;138;142;154mC[38;2;138;142;155mC[38;2;140;142;155mC[38;2;147;149;159mQ[38;2;134;135;140mU[38;2;4;4;6m [38;2;0;0;0m   [38;2;14;12;12m'[38;2;83;79;82mt[38;2;94;92;97mr[38;2;83;82;87mf[38;2;88;86;89mj[38;2;94;92;96mr[38;2;204;202;204mh[38;2;179;180;176mw[38;2;154;158;145mQ[38;2;187;189;174mp[38;2;179;177;168mw[38;2;101;92;91mr[38;2;101;93;96mx[38;2;109;107;113mu[38;2;103;103;112mu[38;2;102;100;110mn[38;2;101;99;110mn[38;2;101;100;112mn[38;2;101;100;113mn[38;2;98;98;111mnn[38;2;101;100;114mn[38;2;103;103;114mu[38;2;102;102;113mn[38;2;103;103;114mu[38;2;101;102;107mn[38;2;111;111;113mv[38;2;150;150;151mL[38;2;185;185;188mp[38;2;158;157;163m0[38;2;103;103;113mu[38;2;127;128;136mY[38;2;100;97;90mr[38;2;78;69;60m?[38;2;83;72;64m?[38;2;86;76;67m1[38;2;87;78;68m1[38;2;90;79;67mt[38;2;91;79;68mt[38;2;95;81;70mt[38;2;97;81;71mf[38;2;99;82;71mf[38;2;99;82;72mf[38;2;100;83;72mff[38;2;102;83;72mf[38;2;103;85;73mj[38;2;105;87;76mj[38;2;105;87;77mj");
  $display("[38;2;169;172;154mZZ[38;2;170;172;155mZ[38;2;169;172;155mZ[38;2;168;172;155mZ[38;2;169;173;156mZ[38;2;161;157;142mQ[38;2;196;184;173mp[38;2;227;211;203mo[38;2;227;210;202mo[38;2;228;208;201mo[38;2;227;208;201mo[38;2;224;208;200ma[38;2;193;181;171mq[38;2;169;161;150mO[38;2;173;171;157mZ[38;2;170;170;156mZ[38;2;168;171;155mOO[38;2;168;171;154mO[38;2;169;171;154mO[38;2;168;171;154mO[38;2;168;171;153mO[38;2;169;172;152mO[38;2;166;168;154mO[38;2;38;39;35ml[38;2;29;9;19m\"[38;2;80;15;48mi[38;2;81;9;49mi[38;2;79;9;48m![38;2;80;10;47m![38;2;81;11;48mi[38;2;82;11;49mi[38;2;85;26;57m+[38;2;202;174;180mp[38;2;228;211;201mo[38;2;223;207;200ma[38;2;224;206;200ma[38;2;225;206;200ma[38;2;226;208;199mo[38;2;229;212;202mo[38;2;202;174;178mp[38;2;108;34;73m?[38;2;118;18;73m?[38;2;114;20;73m?[38;2;112;18;71m-[38;2;107;19;70m-[38;2;109;17;70m-[38;2;110;17;70m--[38;2;112;19;72m-[38;2;111;19;72m-[38;2;107;45;72m1[38;2;159;138;133mC[38;2;171;154;147m0[38;2;125;114;101mv[38;2;83;79;81mt[38;2;88;89;108mr[38;2;201;201;215mh[38;2;245;246;251m@[38;2;248;250;253m@[38;2;252;252;254m$[38;2;239;237;238m8[38;2;184;180;180mq[38;2;250;247;243mB[38;2;255;253;252m$[38;2;252;250;254m$[38;2;244;243;248mB[38;2;208;204;213ma[38;2;145;132;137mJ[38;2;173;154;152m0[38;2;168;149;145mQ[38;2;169;150;146mQ[38;2;170;150;147mQ[38;2;209;190;185mb[38;2;226;207;201mo[38;2;207;188;183mb[38;2;217;198;191mh[38;2;180;163;155mZ[38;2;175;163;158mZ[38;2;213;207;206ma[38;2;225;222;221m#[38;2;233;227;228mW[38;2;235;228;229mW[38;2;238;234;234m&[38;2;232;229;227mW[38;2;218;209;209mo[38;2;171;158;158mO[38;2;149;135;135mJ[38;2;195;180;177mp[38;2;228;211;207m*[38;2;180;164;143mO[38;2;144;135;71mc[38;2;158;148;73mX[38;2;134;108;74mn[38;2;74;21;42m![38;2;83;15;49mi[38;2;99;34;60m-[38;2;102;26;66m-[38;2;101;30;66m-[38;2;107;72;74mf[38;2;109;83;76mj[38;2;108;84;73mj[38;2;108;86;73mj[38;2;112;88;77mr[38;2;115;91;79mr[38;2;114;91;79mr[38;2;115;91;80mr[38;2;115;92;80mr[38;2;114;93;80mr[38;2;113;93;80mr[38;2;111;94;83mx[38;2;106;97;96mx[38;2;104;102;111mn[38;2;98;98;110mn[38;2;97;97;105mx[38;2;99;99;105mn[38;2;103;103;106mn[38;2;105;107;108mu[38;2;106;109;109mu[38;2;111;113;111mv[38;2;119;119;117mc[38;2;43;42;40ml[38;2;40;40;37ml[38;2;47;46;44m![38;2;44;43;43m![38;2;65;61;62m_[38;2;90;87;89mj[38;2;91;89;94mj[38;2;83;82;86mf[38;2;87;85;88mf[38;2;97;95;98mx[38;2;213;211;214mo[38;2;160;160;161mO[38;2;130;133;127mY[38;2;172;173;161mZ[38;2;195;196;184md[38;2;156;155;149mQ[38;2;166;165;161mO[38;2;169;170;166mZ[38;2;175;175;173mw[38;2;174;174;174mw[38;2;168;169;171mZ[38;2;159;161;167mO[38;2;163;166;173mZ[38;2;173;173;181mw[38;2;162;163;170mZ[38;2;147;147;155mL[38;2;145;145;155mL[38;2;148;148;161mQ[38;2;151;151;161mQ[38;2;132;133;135mU[38;2;163;164;156mO[38;2;195;197;183md[38;2;234;236;222mW[38;2;225;226;219m#[38;2;131;132;135mY[38;2;122;121;128mz[38;2;118;110;109mv[38;2;110;94;84mx[38;2;114;95;85mxxx[38;2;114;96;83mxx[38;2;114;96;84mx[38;2;114;95;83mx[38;2;112;94;82mx[38;2;111;93;81mrr[38;2;111;92;80mr[38;2;111;91;80mrrr[38;2;110;92;80mr");
  $display("[38;2;169;172;157mZ[38;2;169;171;156mZ[38;2;170;172;157mZ[38;2;170;172;158mZ[38;2;168;173;157mZ[38;2;171;174;159mZ[38;2;161;154;142mQ[38;2;221;206;197ma[38;2;227;210;202mo[38;2;225;207;200ma[38;2;225;207;199ma[38;2;224;207;199maa[38;2;227;210;202mo[38;2;193;178;169mq[38;2;166;161;147m0[38;2;176;176;160mm[38;2;173;177;159mZ[38;2;172;177;159mZ[38;2;173;176;158mZZZ[38;2;173;175;157mZ[38;2;175;176;157mZ[38;2;167;169;155mO[38;2;38;37;34mI[38;2;51;12;31m;[38;2;83;11;47mi[38;2;80;9;50mii[38;2;80;9;48m![38;2;81;10;48mi[38;2;80;10;47m![38;2;106;50;76m1[38;2;222;196;200ma[38;2;226;208;200mo[38;2;225;206;199ma[38;2;224;207;199maa[38;2;225;208;200mo[38;2;229;213;204m*[38;2;190;162;169mm[38;2;104;29;70m-[38;2;117;19;75m?[38;2;114;20;73m?[38;2;111;18;71m-[38;2;109;18;70m-[38;2;110;17;70m-[38;2;110;17;71m-[38;2;112;18;71m-[38;2;113;20;72m-[38;2;106;18;67m_[38;2;129;76;98mn[38;2;214;197;190mk[38;2;226;211;200mo[38;2;150;143;142mC[38;2;45;52;74m+[38;2;29;42;75mi[38;2;60;66;92m?[38;2;135;135;150mJ[38;2;190;189;198mb[38;2;212;210;216mo[38;2;218;215;222m*[38;2;208;208;213ma[38;2;187;187;192md[38;2;156;159;170mO[38;2;116;123;141mX[38;2;82;91;117mx[38;2;57;68;98m1[38;2;104;101;113mu[38;2;205;189;185mb[38;2;214;195;189mk[38;2;221;202;197ma[38;2;219;200;195mh[38;2;225;206;199ma[38;2;226;207;201mo[38;2;211;192;185mb[38;2;197;178;171mq[38;2;203;186;178md[38;2;198;180;173mp[38;2;206;187;181md[38;2;203;185;179md[38;2;211;194;187mk[38;2;211;196;189mk[38;2;213;198;191mk[38;2;207;193;187mb[38;2;208;191;186mb[38;2;221;203;196ma[38;2;227;209;202mo[38;2;225;206;202mo[38;2;225;208;203mo[38;2;174;159;137m0[38;2;148;138;73mz[38;2;154;140;77mz[38;2;94;54;47m-[38;2;75;12;45m![38;2;85;9;52mi[38;2;105;16;66m_[38;2;116;16;72m-[38;2;100;31;66m-[38;2;114;86;82mr[38;2;114;93;83mx[38;2;112;93;83mx[38;2;111;94;82mr[38;2;112;92;79mr[38;2;112;92;80mr[38;2;112;92;79mr[38;2;112;91;79mrr[38;2;111;91;79mr[38;2;110;91;78mr[38;2;109;92;81mr[38;2;96;85;82mj[38;2;99;98;99mx[38;2;113;113;110mv[38;2;137;138;129mU[38;2;144;146;137mC[38;2;137;141;130mU[38;2;146;150;138mC[38;2;154;157;144mQ[38;2;152;155;140mL[38;2;169;169;153mO[38;2;170;171;156mZ[38;2;143;144;134mJ[38;2;106;106;105mn[38;2;95;93;100mx[38;2;82;80;85mt[38;2;88;86;90mj[38;2;90;89;94mj[38;2;83;82;87mf[38;2;84;83;87mf[38;2;101;99;104mn[38;2;229;227;232mW[38;2;158;157;159m0[38;2;112;112;108mv[38;2;170;171;160mZ[38;2;184;185;170mq[38;2;165;167;152mO[38;2;179;181;166mw[38;2;178;179;162mm[38;2;178;180;162mm[38;2;169;174;162mZ[38;2;106;113;107mu[38;2;91;99;101mx[38;2;124;130;135mY[38;2;167;171;171mZ[38;2;212;215;212mo[38;2;224;226;224mM[38;2;139;139;143mJ[38;2;106;105;115mu[38;2;108;107;117mv[38;2;103;103;107mn[38;2;120;121;117mz[38;2;142;143;136mJ[38;2;146;147;139mC[38;2;132;133;129mY[38;2;102;102;107mn[38;2;125;123;131mX[38;2;120;109;111mv[38;2;107;90;83mr[38;2;111;92;82mrr[38;2;110;91;82mr[38;2;110;92;81mrr[38;2;109;91;80mrr[38;2;108;90;78mrr[38;2;109;91;79mrrrrrr");
  $display("[38;2;207;208;197mh[38;2;206;208;197mh[38;2;208;210;198mh[38;2;209;210;199ma[38;2;206;210;199mh[38;2;209;211;201ma[38;2;183;175;168mw[38;2;214;199;192mk[38;2;226;209;201mo[38;2;224;207;199maaaa[38;2;225;208;200mo[38;2;223;208;198ma[38;2;157;149;136mL[38;2;136;130;116mX[38;2;136;132;117mY[38;2;136;129;115mX[38;2;136;126;114mX[38;2;135;125;112mX[38;2;133;123;111mz[38;2;130;122;110mz[38;2;126;120;107mc[38;2;120;110;103mv[38;2;58;34;41m![38;2;72;12;45m![38;2;82;9;47mi[38;2;77;11;48m![38;2;81;9;49mi[38;2;80;9;49mi[38;2;81;11;48mi[38;2;80;9;46m![38;2;111;56;80mt[38;2;224;201;202ma[38;2;225;207;200ma[38;2;224;207;199maaaa[38;2;230;214;206m*[38;2;181;146;156mO[38;2;104;24;67m-[38;2;118;20;75m?[38;2;114;20;73m?[38;2;111;18;71m-[38;2;110;17;70m--[38;2;110;17;72m-[38;2;113;18;71m-[38;2;114;20;72m-[38;2;102;18;64m_[38;2;159;111;132mU[38;2;232;212;207m*[38;2;219;205;199ma[38;2;99;94;105mx[38;2;70;70;91m1[38;2;91;99;117mn[38;2;38;54;81m+[38;2;31;49;86m+[38;2;31;48;80m~[38;2;35;51;76m~[38;2;43;58;83m_[38;2;43;57;85m_[38;2;34;50;80m~[38;2;28;45;77mii[38;2;28;49;84m~[38;2;32;50;86m+[38;2;130;128;141mU[38;2;228;210;205mo[38;2;226;207;201mo[38;2;225;206;200maa[38;2;225;206;199maa[38;2;226;207;200mo[38;2;196;176;169mq[38;2;212;195;187mk[38;2;194;177;169mq[38;2;224;207;198ma[38;2;225;208;200mo[38;2;223;206;198ma[38;2;224;207;199ma[38;2;226;209;200mo[38;2;226;208;200moo[38;2;224;208;199ma[38;2;224;208;200ma[38;2;225;208;200mo[38;2;224;210;203mo[38;2;163;148;125mC[38;2;155;142;80mX[38;2;137;114;69mu[38;2;76;19;39m![38;2;85;9;52mi[38;2;92;11;53m~[38;2;107;20;69m-[38;2;113;18;70m-[38;2;100;31;68m-[38;2;112;85;81mr[38;2;111;91;79mr[38;2;109;91;79mr[38;2;108;92;79mr[38;2;110;91;77mrrrrr[38;2;111;92;78mrr[38;2;109;92;80mr[38;2;91;81;77mf[38;2;119;118;114mc[38;2;174;176;163mm[38;2;175;177;161mm[38;2;105;107;98mn[38;2;86;89;89mj[38;2;113;116;119mc[38;2;116;118;115mc[38;2;158;160;149mQ[38;2;164;164;154mO[38;2;121;121;118mz[38;2;91;91;92mj[38;2;89;88;92mj[38;2;89;88;94mj[38;2;79;78;83mt[38;2;88;87;92mj[38;2;90;89;94mj[38;2;85;84;89mf[38;2;83;82;87mf[38;2;134;133;138mU[38;2;213;212;217mo[38;2;121;119;123mz[38;2;93;92;90mj[38;2;151;150;143mL[38;2;176;177;164mm[38;2;151;153;138mL[38;2;160;161;146mQ[38;2;172;173;155mZ[38;2;174;175;157mZ[38;2;164;168;158mO[38;2;104;110;104mu[38;2;86;93;92mj[38;2;97;103;104mn[38;2;121;125;121mz[38;2;151;153;147mL[38;2;171;171;169mm[38;2;149;148;152mL[38;2;97;95;106mx[38;2;101;99;112mn[38;2;101;100;107mn[38;2;99;97;106mx[38;2;98;96;105mx[38;2;99;97;106mx[38;2;98;96;106mx[38;2;98;98;106mx[38;2;127;124;132mX[38;2;117;105;108mv[38;2;98;80;74mf[38;2;103;85;75mjj[38;2;101;83;73mf[38;2;102;84;74mf[38;2;101;83;73mfff[38;2;100;82;70mf[38;2;104;86;73mj[38;2;108;90;78mr[38;2;109;91;79mrrrrr");
  $display("[38;2;170;173;156mZ[38;2;172;174;158mZ[38;2;171;174;157mZ[38;2;170;173;157mZ[38;2;170;172;157mZ[38;2;170;174;158mZ[38;2;164;161;147m0[38;2;189;176;166mw[38;2;227;210;202mo[38;2;224;207;199ma[38;2;225;206;199ma[38;2;224;207;199maaa[38;2;228;211;203mo[38;2;191;173;163mw[38;2;106;89;79mj[38;2;109;90;81mrr[38;2;110;89;81mr[38;2;108;88;79mj[38;2;109;88;79mr[38;2;108;88;81mr[38;2;107;89;81mr[38;2;107;77;79mj[38;2;78;25;48mi[38;2;80;9;49mi[38;2;81;9;49mi[38;2;78;10;49m![38;2;80;9;49mi[38;2;79;8;48m![38;2;81;11;48mi[38;2;81;10;46m![38;2;111;59;82mf[38;2;225;201;203ma[38;2;223;208;200ma[38;2;224;207;199ma[38;2;225;207;198maa[38;2;225;206;199ma[38;2;229;212;206m*[38;2;165;125;140mC[38;2;104;21;67m-[38;2;117;19;76m?[38;2;115;20;73m?[38;2;111;18;71m-[38;2;110;17;70m--[38;2;109;18;71m-[38;2;112;18;73m-[38;2;112;18;72m-[38;2;101;19;64m_[38;2;169;124;141mC[38;2;231;214;209m*[38;2;191;175;171mq[38;2;150;138;142mC[38;2;214;201;197mh[38;2;172;164;166mZ[38;2;41;52;82m+[38;2;37;51;91m+[38;2;62;69;97m1[38;2;128;131;151mU[38;2;84;87;112mr[38;2;32;50;85m+[38;2;32;51;89m+[38;2;61;71;95m1[38;2;149;150;159mQ[38;2;106;112;125mv[38;2;43;53;75m+[38;2;140;137;145mJ[38;2;231;214;208m*[38;2;224;207;199maaaa[38;2;225;207;200ma[38;2;225;207;199ma[38;2;217;199;191mh[38;2;203;186;178md[38;2;191;174;166mw[38;2;212;195;187mk[38;2;225;208;200mo[38;2;224;207;199ma[38;2;224;208;200ma[38;2;224;207;199ma[38;2;223;208;199ma[38;2;224;208;199ma[38;2;228;211;202mo[38;2;229;210;201mo[38;2;219;201;193mh[38;2;230;212;211m*[38;2;128;101;103mv[38;2;114;83;61mf[38;2;132;101;72mn[38;2;81;27;42mi[38;2;86;9;52mi[38;2;103;13;63m+[38;2;111;20;70m-[38;2;112;18;72m-[38;2;100;33;67m-[38;2;111;86;79mr[38;2;112;93;79mr[38;2;110;91;78mr[38;2;109;91;78mrrrrr[38;2;109;91;77mr[38;2;110;91;77mrr[38;2;109;92;80mr[38;2;91;81;78mf[38;2;95;91;92mr[38;2;139;137;131mU[38;2;162;164;153m0[38;2;133;135;126mY[38;2;110;113;107mv[38;2;124;127;122mX[38;2;158;162;153m0[38;2;144;147;136mC[38;2;102;102;101mn[38;2;88;87;95mj[38;2;90;90;97mr[38;2;91;90;95mr[38;2;89;87;91mj[38;2;87;87;91mj[38;2;91;90;95mr[38;2;90;90;95mj[38;2;90;89;94mj[38;2;92;91;96mr[38;2;108;106;112mu[38;2;97;96;101mx[38;2;91;89;94mj[38;2;93;92;94mr[38;2;102;101;100mn[38;2;138;138;133mU[38;2;149;147;140mC[38;2;143;141;133mJ[38;2;148;148;138mC[38;2;157;158;147mQQ[38;2;152;154;145mL[38;2;139;143;136mJ[38;2;128;131;126mY[38;2;122;123;121mz[38;2;103;103;104mn[38;2;88;86;93mj[38;2;98;96;105mx[38;2;101;99;110mnn[38;2;100;99;108mn[38;2;101;100;109mn[38;2;101;100;110mnn[38;2;101;100;109mn[38;2;97;98;107mx[38;2;126;124;133mX[38;2;119;108;110mv[38;2;105;87;80mj[38;2;110;91;81mr[38;2;109;91;81mrrrr[38;2;110;92;82mrr[38;2;109;91;80mr[38;2;110;92;81mrr[38;2;110;92;80mr[38;2;109;91;79mrrrr");
  $display("[38;2;217;219;211m*[38;2;216;217;209mo[38;2;216;218;209mo[38;2;217;218;210m*[38;2;220;220;212m*[38;2;219;221;213m*[38;2;223;221;214m*[38;2;200;191;185mb[38;2;212;201;194mh[38;2;224;209;201mo[38;2;225;206;199ma[38;2;224;207;199maaa[38;2;225;208;199ma[38;2;223;205;195ma[38;2;135;117;107mz[38;2;108;90;79mr[38;2;105;86;77mj[38;2;104;84;75mjj[38;2;105;84;76mj[38;2;103;83;75mj[38;2;108;89;79mr[38;2;94;58;65m?[38;2;76;14;47m![38;2;80;9;50mi[38;2;80;8;49m![38;2;80;9;49mii[38;2;80;8;49m![38;2;81;11;48mi[38;2;81;10;47mi[38;2;109;58;81mt[38;2;226;200;203ma[38;2;222;208;200ma[38;2;224;207;199ma[38;2;225;207;198maa[38;2;225;206;200ma[38;2;229;211;206m*[38;2;147;100;120mz[38;2;107;19;69m-[38;2;116;19;77m?[38;2;115;19;73m?[38;2;111;18;71m-[38;2;110;17;70m--[38;2;109;19;71m-[38;2;111;18;75m-[38;2;111;18;74m-[38;2;101;20;64m_[38;2;172;129;143mL[38;2;228;214;204m*[38;2;222;206;194ma[38;2;228;210;205mo[38;2;230;214;204m*[38;2;185;174;173mw[38;2;75;72;92mt[38;2;133;130;143mU[38;2;204;193;193mb[38;2;231;216;207m*[38;2;199;188;182md[38;2;70;75;88m1[38;2;82;85;102mj[38;2;194;187;191md[38;2;234;216;207m*[38;2;227;210;204mo[38;2;175;167;166mZ[38;2;183;173;169mw[38;2;227;211;202mo[38;2;225;209;200mo[38;2;225;209;201mo[38;2;226;210;201mo[38;2;227;211;202mo[38;2;217;201;192mh[38;2;218;202;193mh[38;2;228;212;203mo[38;2;204;188;180md[38;2;210;194;185mb[38;2;229;213;204m*[38;2;228;213;205m*[38;2;228;212;205m*[38;2;229;213;206m*[38;2;229;213;207m*[38;2;227;213;204mo[38;2;220;202;195mh[38;2;194;169;167mw[38;2;132;102;103mv[38;2;148;122;120mY[38;2;220;192;198mh[38;2;102;54;78mt[38;2;74;9;44m![38;2;84;21;54m~[38;2;82;15;52mi[38;2;89;8;55mi[38;2;108;16;68m-[38;2;112;20;69m-[38;2;111;17;74m-[38;2;97;32;64m-[38;2;110;86;77mj[38;2;111;93;78mr[38;2;110;91;77mrr[38;2;109;91;79mrrr[38;2;109;91;78mr[38;2;109;91;77mr[38;2;110;92;77mr[38;2;110;92;78mr[38;2;110;91;78mr[38;2;95;83;83mj[38;2;96;91;101mx[38;2;69;66;73m?[38;2;80;79;82mt[38;2;96;96;98mx[38;2;100;100;102mxx[38;2;92;93;95mr[38;2;83;82;87mf[38;2;82;80;87mf[38;2;84;81;85mf[38;2;83;80;82mt[38;2;83;79;80mt[38;2;84;78;77mt[38;2;84;78;79mt[38;2;83;77;78mt[38;2;83;77;79mt[38;2;84;76;77mt[38;2;87;76;75mt[38;2;85;74;73m1[38;2;84;73;72m1[38;2;85;75;74mt[38;2;83;74;73m1[38;2;80;71;68m?[38;2;78;70;65m?[38;2;80;70;70m?[38;2;77;69;71m?[38;2;74;71;73m?[38;2;72;71;74m?[38;2;71;69;72m?[38;2;68;67;71m-[38;2;69;69;75m?[38;2;76;77;83mt[38;2;88;87;94mj[38;2;97;96;104mx[38;2;101;100;109mn[38;2;101;99;111mnn[38;2;101;99;112mn[38;2;101;100;111mn[38;2;101;101;109mn[38;2;100;101;108mn[38;2;101;101;109mn[38;2;101;101;108mn[38;2;97;100;109mn[38;2;126;125;136mY[38;2;120;110;110mv[38;2;106;89;81mr[38;2;107;89;79mj[38;2;106;88;78mj[38;2;107;89;79mj[38;2;106;88;78mjjjjjjj[38;2;105;87;76mj[38;2;104;86;74mj[38;2;106;88;76mj[38;2;110;92;80mr[38;2;109;91;79mr");
  $display("[38;2;239;239;236m8[38;2;238;238;234m&[38;2;238;239;235m&[38;2;239;240;236m8[38;2;241;241;237m8[38;2;240;241;237m8[38;2;243;242;238m8[38;2;237;234;231m&[38;2;196;189;185md[38;2;223;209;202mo[38;2;226;207;198ma[38;2;224;207;199maaaa[38;2;230;212;203m*[38;2;182;163;155mZ[38;2;103;85;76mj[38;2;107;88;79mj[38;2;106;87;78mjj[38;2;106;87;77mj[38;2;105;89;79mj[38;2;110;87;84mr[38;2;80;35;52m+[38;2;78;11;50mi[38;2;81;9;50mi[38;2;80;8;48m!![38;2;79;8;48m![38;2;79;10;49mi[38;2;81;11;48mi[38;2;79;11;47m![38;2;103;51;74m1[38;2;225;196;199ma[38;2;224;209;201mo[38;2;223;208;200ma[38;2;226;208;200mo[38;2;226;209;201mo[38;2;226;209;203mo[38;2;221;197;197mh[38;2;121;63;88mj[38;2;114;19;70m-[38;2;115;19;76m?[38;2;114;19;73m-[38;2;111;17;70m-[38;2;111;17;69m--[38;2;110;18;72m-[38;2;113;17;74m--[38;2;102;17;67m_[38;2;174;126;150mL[38;2;235;217;214m#[38;2;227;209;201mo[38;2;227;208;203mo[38;2;216;197;190mk[38;2;156;135;133mJ[38;2;190;172;175mq[38;2;228;212;209m*[38;2;233;215;208m*[38;2;232;213;206m*[38;2;233;215;209m*[38;2;205;192;185mb[38;2;212;199;192mk[38;2;232;215;209m*[38;2;231;211;204m*[38;2;230;212;203m*[38;2;230;212;204m*[38;2;228;207;202mo[38;2;221;200;197ma[38;2;217;196;193mh[38;2;214;192;189mk[38;2;210;187;184mb[38;2;205;182;180md[38;2;195;171;170mw[38;2;190;166;165mm[38;2;189;165;163mm[38;2;179;153;151mO[38;2;184;156;155mZ[38;2;180;151;150mO[38;2;177;147;148m0[38;2;173;141;145mQ[38;2;168;135;139mL[38;2;158;124;129mU[38;2;134;101;106mv[38;2;112;86;91mx[38;2;135;112;121mz[38;2;116;86;100mx[38;2;92;51;68m?[38;2;94;48;69m?[38;2;75;16;47mi[38;2;83;11;52mi[38;2;81;9;52mi[38;2;81;8;53mi[38;2;92;11;60m~[38;2;108;18;70m-[38;2;111;20;70m-[38;2;111;17;74m-[38;2;98;31;65m-[38;2;111;86;77mj[38;2;110;93;78mr[38;2;110;93;80mr[38;2;111;92;81mr[38;2;111;93;80mr[38;2;111;93;81mr[38;2;111;93;82mr[38;2;111;93;81mr[38;2;110;92;81mr[38;2;111;93;80mr[38;2;111;93;79mr[38;2;113;93;81mr[38;2;88;75;74mt[38;2;71;67;76m?[38;2;61;60;69m_[38;2;57;56;62m+[38;2;60;59;65m__[38;2;59;58;63m__[38;2;61;58;67m_[38;2;60;54;59m+[38;2;68;57;55m_[38;2;75;59;53m_[38;2;75;58;50m__[38;2;76;58;51m__[38;2;77;58;52m_[38;2;77;58;51m___[38;2;76;58;51m_[38;2;77;58;51m_[38;2;78;60;52m_[38;2;78;61;52m_[38;2;78;60;51m_[38;2;77;60;55m-[38;2;66;52;53m+[38;2;64;57;61m_[38;2;60;59;63m_[38;2;62;61;67m_[38;2;73;72;78m1[38;2;82;81;88mf[38;2;86;85;93mj[38;2;86;84;94mj[38;2;81;80;89mf[38;2;81;80;88mf[38;2;81;80;89mf[38;2;81;80;90mf[38;2;80;78;89mt[38;2;78;77;87mt[38;2;78;78;86mt[38;2;77;77;85mtt[38;2;78;77;85mt[38;2;72;75;83m1[38;2;112;111;120mv[38;2;122;111;113mc[38;2;104;87;80mj[38;2;106;88;78mjj[38;2;105;87;77mjjjj[38;2;108;90;80mr[38;2;109;91;81mrr[38;2;109;91;82mr[38;2;110;92;81mr[38;2;108;90;78mr[38;2;109;91;79mrrr");
  $display("[38;2;178;180;167mw[38;2;177;179;166mw[38;2;178;180;166mw[38;2;178;180;167mwwww[38;2;188;190;178mp[38;2;193;190;180mp[38;2;208;197;187mk[38;2;226;209;201mo[38;2;225;208;200mo[38;2;226;209;201mooo[38;2;228;209;202mo[38;2;218;198;192mh[38;2;125;106;99mv[38;2;110;91;83mr[38;2;111;93;82mr[38;2;110;92;82mrr[38;2;109;93;83mr[38;2;106;77;79mj[38;2;75;23;46mi[38;2;80;11;49mi[38;2;80;9;49miii[38;2;79;9;49m![38;2;79;10;49mi[38;2;81;11;48mi[38;2;77;11;46m![38;2;105;57;79mt[38;2;224;199;201ma[38;2;199;186;177mp[38;2;181;165;157mZ[38;2;183;165;157mZ[38;2;207;192;184mb[38;2;229;212;207m*[38;2;193;163;168mw[38;2;99;30;66m-[38;2;115;20;74m?[38;2;113;20;75m?[38;2;113;18;72m-[38;2;111;16;71m-[38;2;111;17;71m---[38;2;114;17;72m--[38;2;107;19;70m-[38;2;120;64;90mj[38;2;183;152;155mO[38;2;220;190;190mk[38;2;231;210;211m*[38;2;212;187;189mb[38;2;84;48;55m_[38;2;96;55;65m?[38;2;122;83;92mx[38;2;140;102;110mc[38;2;152;115;123mY[38;2;158;119;128mU[38;2;160;121;128mU[38;2;153;115;123mY[38;2;144;106;116mz[38;2;136;98;110mv[38;2;130;92;104mu[38;2;123;85;97mn[38;2;119;81;93mx[38;2;114;76;87mr[38;2;111;73;83mj[38;2;109;72;81mj[38;2;113;76;86mj[38;2;114;78;89mr[38;2;117;83;94mx[38;2;120;88;98mn[38;2;123;92;102mn[38;2;116;85;95mx[38;2;131;101;111mv[38;2;138;110;119mz[38;2;141;114;123mX[38;2;146;119;129mY[38;2;150;125;135mU[38;2;140;116;125mX[38;2;185;169;175mw[38;2;223;218;220m#[38;2;229;221;224mM[38;2;123;101;108mv[38;2;88;51;62m-[38;2;139;95;114mc[38;2;79;20;52mi[38;2;80;10;50mi[38;2;81;10;51mi[38;2;85;10;54mi[38;2;102;15;66m_[38;2;111;17;71m-[38;2;112;19;71m-[38;2;114;17;76m?[38;2;99;29;64m-[38;2;103;75;71mf[38;2;101;83;73mf[38;2;100;83;74mf[38;2;100;82;71mf[38;2;98;80;67mt[38;2;97;79;66mt[38;2;93;75;64m1[38;2;91;72;64m1[38;2;90;71;64m1[38;2;90;72;63m1[38;2;92;74;62m1[38;2;94;74;63m1[38;2;74;62;58m-[38;2;60;57;60m+[38;2;61;60;66m__[38;2;60;59;65m_[38;2;59;58;64m_[38;2;60;59;64m_[38;2;61;60;65m_[38;2;61;59;66m_[38;2;60;53;57m+[38;2;69;55;54m+[38;2;78;60;52m_[38;2;80;59;49m_[38;2;78;59;51m_[38;2;77;58;50m_[38;2;78;57;50m_[38;2;79;58;51m_[38;2;78;58;51m_[38;2;77;58;51m__[38;2;78;59;52m_[38;2;77;58;50m_[38;2;78;60;50m_[38;2;79;61;51m__[38;2;80;62;55m-[38;2;67;53;54m+[38;2;63;57;63m_[38;2;61;61;64m_[38;2;61;61;67m_[38;2;62;61;67m_[38;2;61;60;66m_[38;2;60;59;65m_[38;2;60;59;64m_[38;2;59;58;64m_[38;2;60;59;64m__[38;2;59;59;64m_[38;2;60;59;64m_[38;2;59;58;64m_[38;2;55;54;59m+[38;2;57;55;61m+[38;2;57;56;62m+[38;2;58;57;63m+[38;2;54;56;64m+[38;2;106;105;112mu[38;2;122;112;114mc[38;2;106;89;83mr[38;2;110;92;82mr[38;2;108;90;80mr[38;2;107;89;79mj[38;2;106;88;78mjj[38;2;107;88;78mj[38;2;110;92;82mr[38;2;110;92;80mrr[38;2;109;92;80mrr[38;2;109;91;79mrrrr");
  $display("[38;2;155;157;145mQ[38;2;155;157;146mQ[38;2;154;155;144mQ[38;2;153;155;143mL[38;2;153;155;144mL[38;2;153;155;143mL[38;2;150;152;141mL[38;2;147;149;136mC[38;2;149;149;136mC[38;2;148;140;130mJ[38;2;220;205;197ma[38;2;214;196;189mk[38;2;206;189;181mb[38;2;205;188;180md[38;2;204;187;179md[38;2;214;196;188mk[38;2;230;212;204m*[38;2;172;154;147m0[38;2;105;87;78mj[38;2;112;94;83mx[38;2;111;93;83mr[38;2;110;93;82mr[38;2;111;92;83mr[38;2;99;71;72mt[38;2;73;18;42m![38;2;80;10;48mi[38;2;79;9;49m!!![38;2;79;10;49mi[38;2;78;9;48m![38;2;82;11;50mi[38;2;75;11;45m![38;2;146;105;122mX[38;2;232;212;211m*[38;2;215;204;195mh[38;2;217;199;193mh[38;2;214;197;191mk[38;2;217;202;193mh[38;2;230;213;206m*[38;2;172;143;149mQ[38;2;92;21;61m+[38;2;112;22;75m?[38;2;111;21;75m?[38;2;112;17;73m-[38;2;111;17;74m-[38;2;111;18;74m-[38;2;106;14;69m_[38;2;109;18;70m-[38;2;114;18;71m-[38;2;114;18;72m-[38;2;107;20;69m-[38;2;117;62;87mj[38;2;100;63;71mt[38;2;92;47;59m-[38;2;122;77;94mx[38;2;135;92;106mv[38;2;82;36;52m+[38;2;130;96;111mv[38;2;194;180;185mp[38;2;176;163;166mZ[38;2;166;150;154m0[38;2;164;145;150mQ[38;2;164;143;149mQ[38;2;165;146;153mQ[38;2;145;129;135mU[38;2;183;169;175mw[38;2;194;182;187mp[38;2;203;193;197mk[38;2;209;201;204mh[38;2;216;208;212mo[38;2;216;209;212mo[38;2;198;193;195mb[38;2;238;234;236m&[38;2;242;237;240m8[38;2;247;243;246mB[38;2;252;248;251m@[38;2;254;252;255m$[38;2;213;215;216mo[38;2;253;253;255m$[38;2;255;255;255m$$$$[38;2;218;214;216m*[38;2;255;255;255m$$[38;2;208;201;202mh[38;2;95;69;75mt[38;2;179;150;154mO[38;2;188;154;167mZ[38;2;70;15;46m![38;2;81;10;51mi[38;2;81;9;51mi[38;2;92;11;57m~[38;2;110;17;69m-[38;2;113;15;71m-[38;2;112;18;70m-[38;2;115;16;76m?[38;2;98;24;64m_[38;2;81;51;54m_[38;2;77;59;51m_[38;2;77;60;50m_[38;2;79;60;51m_[38;2;79;61;49m_[38;2;78;60;49m_[38;2;78;60;50m_[38;2;77;59;51m_[38;2;75;57;49m_[38;2;74;55;47m+[38;2;77;59;49m_[38;2;81;62;50m-[38;2;67;55;50m+[38;2;61;58;60m+[38;2;60;59;64m_[38;2;61;60;65m_[38;2;72;72;77m?[38;2;77;76;81mt[38;2;65;64;68m-[38;2;59;58;63m_[38;2;62;60;67m_[38;2;62;54;59m+[38;2;70;56;55m_[38;2;79;61;54m-[38;2;80;62;51m-[38;2;79;60;53m-[38;2;75;56;48m+[38;2;74;55;47m+[38;2;75;56;49m_[38;2;74;56;49m+[38;2;74;55;48m++[38;2;75;56;49m_[38;2;75;57;49m_[38;2;74;56;46m++[38;2;77;59;49m_[38;2;77;61;54m-[38;2;64;54;54m+[38;2;61;57;62m_[38;2;59;61;64m_[38;2;61;60;65m__[38;2;60;59;64m_[38;2;60;59;65m_[38;2;61;60;64m_[38;2;61;60;65m_[38;2;61;60;64m___[38;2;60;59;64m_[38;2;69;69;73m?[38;2;147;147;150mL[38;2;202;202;204mh[38;2;161;161;164mO[38;2;87;86;90mj[38;2;55;56;64m+[38;2;110;108;116mv[38;2;122;111;114mc[38;2;106;88;83mr[38;2;109;91;81mr[38;2;109;92;82mr[38;2;110;93;83mrrrrr[38;2;110;91;79mrrrr[38;2;111;92;80mrrr[38;2;110;91;80mr");
  $display("[38;2;93;92;95mrr[38;2;92;92;94mr[38;2;91;91;93mj[38;2;92;91;94mrr[38;2;91;91;93mjj[38;2;93;90;90mj[38;2;80;70;69m?[38;2;188;171;169mw[38;2;216;198;191mk[38;2;189;172;164mww[38;2;199;183;174mp[38;2;217;200;192mh[38;2;226;209;201mo[38;2;221;204;196ma[38;2;125;107;99mv[38;2;88;70;60m?[38;2;92;74;64m11[38;2;91;72;63m1[38;2;81;55;55m_[38;2;73;15;41m![38;2;79;10;48m![38;2;80;9;49miii[38;2;80;9;48m![38;2;79;11;48mi[38;2;83;11;52mi[38;2;75;14;47m![38;2;174;140;151mQ[38;2;232;212;208m*[38;2;222;208;199ma[38;2;223;208;202mo[38;2;224;209;202mo[38;2;224;208;199ma[38;2;230;214;206m*[38;2;161;134;141mC[38;2;87;19;56m~[38;2;110;21;73m-[38;2;111;20;74m-[38;2;114;17;73m-[38;2;113;18;74m-[38;2;109;19;72m-[38;2;97;11;61m+[38;2;104;16;67m_[38;2;111;17;70m-[38;2;113;17;71m-[38;2;105;17;67m_[38;2;139;86;110mv[38;2;209;186;188mb[38;2;156;125;129mU[38;2;96;52;67m?[38;2;75;25;42mi[38;2;81;28;48m~[38;2;119;85;101mn[38;2;208;203;207ma[38;2;254;255;254m$[38;2;254;254;254m$[38;2;255;255;255m$$$[38;2;217;219;218m*[38;2;242;245;244mB[38;2;255;255;255m$[38;2;254;255;255m$[38;2;254;254;254m$[38;2;251;249;250m@[38;2;247;245;246mB[38;2;205;202;203mh[38;2;225;222;223m#[38;2;219;215;217m*[38;2;206;201;202mh[38;2;191;183;186mp[38;2;176;167;170mm[38;2;143;132;136mU[38;2;157;145;150mL[38;2;157;143;148mL[38;2;151;136;141mC[38;2;143;128;133mU[38;2;135;121;123mX[38;2;116;102;102mu[38;2;127;114;115mc[38;2;125;113;113mc[38;2;104;83;87mj[38;2;78;48;54m_[38;2;203;179;182md[38;2;158;124;136mJ[38;2;68;10;41ml[38;2;84;10;52mi[38;2;83;9;52mi[38;2;97;13;60m+[38;2;112;18;70m-[38;2;114;15;71m-[38;2;110;18;69m-[38;2;112;16;75m-[38;2;98;23;65m_[38;2;81;50;54m_[38;2;79;61;52m-[38;2;78;61;50m_[38;2;80;60;53m-[38;2;80;62;52m----[38;2;81;63;53m-[38;2;79;61;51m__[38;2;81;61;51m-[38;2;69;55;52m+[38;2;59;56;60m+[38;2;61;60;66m_[38;2;105;105;105mn[38;2;134;134;134mU[38;2;219;219;218m*[38;2;201;200;201mk[38;2;82;80;86mt[38;2;59;57;64m_[38;2;62;55;59m+[38;2;72;57;56m_[38;2;78;61;53m-[38;2;79;61;50m_[38;2;81;61;53m-[38;2;79;59;50m_[38;2;77;59;50m_[38;2;76;59;52m_[38;2;75;59;52m_[38;2;78;59;52m_[38;2;77;58;51m_[38;2;78;59;52m_[38;2;78;59;51m_[38;2;78;61;50m__[38;2;79;61;51m_[38;2;78;61;55m-[38;2;67;53;55m+[38;2;64;58;63m_[38;2;61;60;64m_[38;2;61;60;65m__[38;2;59;58;63m__[38;2;60;58;64m_[38;2;60;59;64m_[38;2;61;60;65m___[38;2;58;57;62m+[38;2;94;93;98mr[38;2;141;141;143mJ[38;2;144;144;146mC[38;2;119;119;120mz[38;2;98;98;101mx[38;2;57;58;66m_[38;2;112;109;117mv[38;2;125;113;116mc[38;2;107;89;83mr[38;2;111;91;82mrr[38;2;110;91;82mr[38;2;109;90;81mr[38;2;108;89;79mr[38;2;107;88;78mj[38;2;106;86;77mj[38;2;105;85;74mj[38;2;103;83;72mff[38;2;102;82;71mf[38;2;100;80;69mf[38;2;99;79;68mt[38;2;98;78;67mt[38;2;97;77;66mt");
  $display("[38;2;89;88;94mjjjjjjj[38;2;90;89;94mj[38;2;93;90;94mr[38;2;74;64;64m-[38;2;126;111;104mv[38;2;232;214;206m*[38;2;230;212;204m*[38;2;228;210;203mo[38;2;227;209;202mo[38;2;225;208;200mo[38;2;224;207;199ma[38;2;228;211;203mo[38;2;199;181;173mp[38;2;91;72;64m1[38;2;79;61;52m-[38;2;81;63;54m-[38;2;80;62;53m-[38;2;80;54;53m_[38;2;73;20;42m![38;2;81;11;50mi[38;2;80;9;50mi[38;2;80;9;49mii[38;2;79;9;47m![38;2;78;12;48mi[38;2;83;10;51mi[38;2;84;23;55m~[38;2;195;166;173mw[38;2;230;210;204mo[38;2;225;207;197ma[38;2;223;207;198ma[38;2;223;208;200ma[38;2;223;208;198ma[38;2;232;214;207m*[38;2;160;130;138mC[38;2;83;17;53m~[38;2;110;20;71m-[38;2;111;20;73m-[38;2;114;18;72m-[38;2;113;19;72m-[38;2;106;18;68m-[38;2;89;8;54mi[38;2;99;13;62m+[38;2;111;17;70m-[38;2;113;18;72m-[38;2;107;18;69m-[38;2;121;65;90mr[38;2;201;180;177mp[38;2;236;215;208m*[38;2;219;194;194mh[38;2;163;137;143mL[38;2;98;57;73m1[38;2;91;52;70m?[38;2;193;181;189mp[38;2;240;237;241m8[38;2;252;250;253m@[38;2;243;239;242m8[38;2;232;228;229mW[38;2;218;213;214m*[38;2;184;177;179mq[38;2;158;149;150mQ[38;2;163;154;155m0[38;2;146;135;138mJ[38;2;131;117;123mz[38;2;116;99;106mu[38;2;101;85;90mr[38;2;81;66;70m?[38;2;76;57;62m-[38;2;71;48;56m+[38;2;64;43;49m~[38;2;60;38;43mi[38;2;59;34;39m![38;2;60;34;39m![38;2;60;32;38m!![38;2;57;32;37m![38;2;57;32;36ml[38;2;58;32;36m![38;2;60;35;38m![38;2;58;34;36m![38;2;60;33;36m![38;2;63;29;35m![38;2;87;52;58m-[38;2;215;194;194mk[38;2;133;96;111mv[38;2;71;8;42ml[38;2;84;11;52mi[38;2;84;9;51mi[38;2;96;12;59m+[38;2;112;16;69m-[38;2;113;16;71m-[38;2;109;18;69m-[38;2;114;15;75m-[38;2;101;22;66m_[38;2;82;49;55m_[38;2;80;61;53m-[38;2;78;61;50m_[38;2;80;60;52m-[38;2;80;62;52m---[38;2;80;62;51m-[38;2;79;61;50m__[38;2;79;61;51m_[38;2;81;61;51m-[38;2;69;56;53m+[38;2;60;57;61m+[38;2;62;61;66m_[38;2;84;84;88mf[38;2;90;89;94mj[38;2;120;119;124mz[38;2;144;143;147mC[38;2;87;86;92mj[38;2;59;57;65m_[38;2;62;55;60m+[38;2;72;57;56m_[38;2;78;61;53m-[38;2;79;61;50m_[38;2;81;61;53m-[38;2;80;61;52m-[38;2;80;62;52m-[38;2;79;62;53m-[38;2;79;62;54m-[38;2;80;61;53m--[38;2;80;62;53m--[38;2;81;62;52m---[38;2;80;61;54m-[38;2;68;54;54m+[38;2;65;57;64m_[38;2;62;60;65m_[38;2;61;60;65m__[38;2;60;59;64m____[38;2;61;60;65m____[38;2;60;59;64m_[38;2;67;67;70m-[38;2;71;71;74m?[38;2;72;71;75m?[38;2;62;61;65m_[38;2;56;57;64m+[38;2;109;107;116mv[38;2;117;107;109mv[38;2;83;64;58m-[38;2;89;67;59m??[38;2;88;66;58m?[38;2;87;65;57m?[38;2;85;63;55m-[38;2;84;62;54m-[38;2;83;62;53m-[38;2;81;61;51m----[38;2;80;60;50m____");
  $display("[38;2;89;88;93mjjjjjjj[38;2;90;89;93mj[38;2;93;89;94mr[38;2;78;67;68m?[38;2;81;65;57m-[38;2;192;173;165mw[38;2;232;213;206m*[38;2;226;207;200moo[38;2;224;207;199maaa[38;2;230;212;205m*[38;2;164;145;138mL[38;2;79;60;53m-[38;2;83;64;57m-[38;2;81;64;54m-[38;2;82;59;53m-[38;2;73;29;44mi[38;2;77;11;48m![38;2;80;9;49miii[38;2;79;9;48m![38;2;78;11;49mi[38;2;83;9;49mi[38;2;100;42;70m?[38;2;216;192;194mk[38;2;225;210;202mo[38;2;224;207;198ma[38;2;224;207;197ma[38;2;224;207;198ma[38;2;222;208;197ma[38;2;232;213;208m*[38;2;156;123;132mU[38;2;80;14;49mi[38;2;106;17;67m_[38;2;111;19;71m-[38;2;113;16;71m-[38;2;109;18;71m-[38;2;102;16;66m_[38;2;87;7;53mi[38;2;95;10;56m~[38;2;110;18;68m-[38;2;114;19;72m-[38;2;109;18;71m-[38;2;114;53;83mf[38;2;174;153;150m0[38;2;225;206;195ma[38;2;229;210;203mo[38;2;234;219;213m#[38;2;161;132;137mC[38;2;75;32;47m~[38;2;138;110;122mz[38;2;135;117;125mX[38;2;116;102;106mu[38;2;94;76;80mf[38;2;79;60;63m-[38;2;69;48;52m+[38;2;62;40;45mi[38;2;57;35;39m![38;2;53;33;34ml[38;2;55;31;35ml[38;2;61;34;39m![38;2;69;37;42mi[38;2;76;41;46m~[38;2;79;42;48m+[38;2;81;42;49m+[38;2;80;43;48m+[38;2;75;41;46m~[38;2;69;37;42mi[38;2;66;35;38mi[38;2;63;35;36m![38;2;63;37;38mi[38;2;63;37;40mi[38;2;62;36;40mi[38;2;62;37;40mi[38;2;61;37;39m![38;2;61;36;39m![38;2;61;37;39m![38;2;63;36;39mi[38;2;62;29;34ml[38;2;111;74;80mj[38;2;229;200;201ma[38;2;113;69;87mj[38;2;73;9;45m![38;2;85;10;51mi[38;2;84;9;50mi[38;2;97;11;58m+[38;2;112;15;67m-[38;2;113;15;71m-[38;2;110;18;69m-[38;2;115;16;75m-[38;2;102;21;66m_[38;2;84;47;55m_[38;2;81;61;54m-[38;2;78;62;49m_[38;2;80;61;51m-[38;2;80;62;52m---[38;2;80;62;50m-[38;2;79;61;48m_[38;2;78;60;49m_[38;2;79;61;51m_[38;2;81;61;52m-[38;2;69;56;53m+[38;2;60;58;62m_[38;2;61;60;64m_[38;2;60;59;64m_[38;2;66;65;70m-[38;2;64;63;68m-[38;2;67;65;70m-[38;2;60;59;66m_[38;2;62;60;68m_[38;2;61;53;60m+[38;2;69;55;55m+[38;2;79;62;54m-[38;2;80;62;51m-[38;2;81;61;54m-[38;2;80;62;52m--------[38;2;81;61;52m---[38;2;79;62;54m-[38;2;68;56;55m+[38;2;63;57;64m_[38;2;61;59;65m_[38;2;61;60;65m___________[38;2;60;59;64m_[38;2;59;58;63m_[38;2;60;59;64m__[38;2;56;56;63m+[38;2;106;105;115mu[38;2;114;105;107mu[38;2;74;57;49m_[38;2;80;60;51m_[38;2;81;61;52m--------------");
  $display("[38;2;89;88;93mjjjjjjj[38;2;89;89;93mj[38;2;91;88;93mj[38;2;78;69;70m?[38;2;76;61;53m_[38;2;126;107;99mv[38;2;227;208;201mo[38;2;226;208;200mo[38;2;225;206;199ma[38;2;224;207;199maaa[38;2;225;208;200mo[38;2;225;207;199ma[38;2;119;100;93mn[38;2;77;59;51m_[38;2;81;62;52m-[38;2;82;61;53m-[38;2;80;44;51m+[38;2;71;14;42m![38;2;80;9;49miii[38;2;80;9;48m![38;2;81;10;51mi[38;2;80;8;48m![38;2;117;66;88mj[38;2;226;205;203mo[38;2;223;208;200ma[38;2;223;208;198maa[38;2;224;207;198ma[38;2;221;208;197ma[38;2;231;212;208m*[38;2;151;114;127mY[38;2;81;12;49mi[38;2;98;15;61m+[38;2;109;18;69m-[38;2;115;15;70m-[38;2;110;18;71m-[38;2;99;13;62m+[38;2;86;6;51mi[38;2;90;7;53mi[38;2;109;17;69m-[38;2;115;19;73m?[38;2;111;18;73m-[38;2;104;39;73m?[38;2;158;131;133mJ[38;2;201;186;173mp[38;2;227;210;199mo[38;2;227;213;204mo[38;2;191;170;165mw[38;2;82;40;53m+[38;2;69;28;44mi[38;2;60;29;38m![38;2;59;32;39m![38;2;62;35;40m![38;2;64;36;41mi[38;2;62;36;39m![38;2;66;35;38mi[38;2;86;44;49m+[38;2;115;56;65mt[38;2;142;69;81mx[38;2;163;78;93mv[38;2;175;84;97mc[38;2;183;85;99mz[38;2;187;86;101mX[38;2;185;87;101mX[38;2;182;86;98mz[38;2;179;84;96mz[38;2;168;79;91mv[38;2;150;71;81mx[38;2;121;56;64mt[38;2;93;39;45m+[38;2;68;34;35m![38;2;59;37;35m![38;2;61;37;38m![38;2;63;35;39m![38;2;62;36;38m![38;2;59;37;38m![38;2;61;36;39m![38;2;59;28;33ml[38;2;128;94;99mu[38;2;228;193;197ma[38;2;95;44;66m-[38;2;76;10;46m![38;2;83;11;51mi[38;2;83;8;49mi[38;2;94;10;56m~[38;2;111;17;67m-[38;2;114;15;70m-[38;2;111;17;67m-[38;2;113;16;74m-[38;2;99;23;66m_[38;2;82;47;53m_[38;2;80;60;51m_[38;2;79;62;49m_[38;2;80;61;51m-[38;2;80;62;51m-[38;2;79;61;51m_[38;2;77;59;50m_[38;2;77;59;48m_[38;2;76;58;47m__[38;2;77;59;49m_[38;2;78;59;49m_[38;2;67;55;51m+[38;2;61;57;60m+[38;2;61;60;64m_[38;2;61;60;65m_[38;2;60;59;64m_[38;2;59;58;63m_[38;2;60;59;64m_[38;2;60;60;67m_[38;2;61;60;68m_[38;2;61;53;60m+[38;2;70;55;54m+[38;2;80;61;54m-[38;2;80;62;51m-[38;2;81;61;54m-[38;2;80;62;52m--------[38;2;81;61;52m---[38;2;79;62;53m-[38;2;66;54;53m+[38;2;62;56;63m_[38;2;61;59;66m_[38;2;61;60;66m_[38;2;61;60;65m_[38;2;60;59;64m_[38;2;61;60;65m_______[38;2;61;60;66m__[38;2;61;60;65m___[38;2;56;56;64m+[38;2;100;100;111mn[38;2;113;105;107mu[38;2;74;58;51m_[38;2;79;61;51m_[38;2;79;61;52m--[38;2;79;61;51m_[38;2;79;60;50m_[38;2;78;59;50m____[38;2;79;60;50m_[38;2;79;60;51m_[38;2;79;59;50m___[38;2;78;58;50m_");
  $display("[38;2;89;88;93mjjjjjjj[38;2;88;87;91mj[38;2;88;87;92mj[38;2;76;70;70m?[38;2;80;65;57m-[38;2;83;65;57m-[38;2;184;167;159mm[38;2;229;212;204m*[38;2;224;207;199maaaaa[38;2;230;213;205m*[38;2;189;172;164mw[38;2;80;63;55m-[38;2;79;59;51m_[38;2;78;61;52m_[38;2;81;57;55m-[38;2;72;28;44mi[38;2;74;11;46m![38;2;80;9;48m![38;2;81;8;49mi[38;2;79;9;49m![38;2;82;9;50mi[38;2;77;8;48m![38;2;137;97;114mc[38;2;230;211;206m*[38;2;225;208;199ma[38;2;224;207;199maa[38;2;225;207;198ma[38;2;222;208;197ma[38;2;231;210;208m*[38;2;139;98;114mc[38;2;78;10;46m![38;2;89;11;53m~[38;2;103;17;67m_[38;2;114;16;70m-[38;2;110;18;70m-[38;2;95;11;58m~[38;2;83;7;49mi[38;2;87;8;51mi[38;2;106;18;66m_[38;2;112;19;71m-[38;2;110;20;71m-[38;2;101;28;65m-[38;2;150;113;122mY[38;2;176;159;150mO[38;2;223;205;194ma[38;2;227;209;201mo[38;2;217;197;193mh[38;2;97;60;74m1[38;2;75;30;48m~[38;2;68;33;44mi[38;2;64;37;41mi[38;2;66;33;37m![38;2;72;34;38mi[38;2;104;49;56m?[38;2;150;70;82mx[38;2;184;86;100mz[38;2;194;91;103mY[38;2;198;94;107mU[38;2;200;96;109mU[38;2;200;96;110mU[38;2;202;98;112mU[38;2;204;100;115mJ[38;2;205;102;116mJ[38;2;207;100;115mJ[38;2;208;101;116mJ[38;2;207;100;114mJ[38;2;204;98;112mJ[38;2;201;96;108mU[38;2;189;88;101mX[38;2;153;73;81mn[38;2;100;49;48m-[38;2;66;33;33m![38;2;62;34;39m![38;2;63;36;39mi[38;2;62;36;37m![38;2;63;36;38m![38;2;59;29;34ml[38;2;152;121;128mU[38;2;215;180;188mb[38;2;80;27;52m~[38;2;81;10;50mi[38;2;83;10;52mi[38;2;79;9;48m![38;2;88;8;53mi[38;2;106;15;65m_[38;2;110;13;68m_[38;2;110;18;68m-[38;2;112;16;72m-[38;2;98;23;63m_[38;2;81;48;51m_[38;2;79;60;49m_[38;2;80;62;48m_[38;2;81;60;52m-[38;2;79;61;49m_[38;2;79;61;50m_[38;2;75;57;49m_[38;2;75;56;48m+[38;2;76;58;48m_[38;2;78;60;50m_[38;2;79;61;51m_[38;2;78;62;50m_[38;2;66;54;50m+[38;2;63;57;60m_[38;2;61;60;63m_[38;2;61;60;65m___[38;2;59;58;63m_[38;2;60;60;66m_[38;2;61;60;68m_[38;2;60;53;60m+[38;2;72;55;55m_[38;2;81;60;54m-[38;2;81;61;51m-[38;2;81;61;54m-[38;2;80;62;52m--------[38;2;81;61;52m---[38;2;79;63;52m-[38;2;66;54;53m+[38;2;62;56;63m_[38;2;61;60;68m__[38;2;61;60;66m_[38;2;61;60;65m_[38;2;61;60;64m_[38;2;61;60;65m___[38;2;61;60;64m_[38;2;61;60;65m_[38;2;61;60;66m_[38;2;61;60;68m__[38;2;61;60;66m_[38;2;61;60;65m_[38;2;61;60;64m_[38;2;56;56;65m+[38;2;95;97;109mx[38;2;113;105;109mu[38;2;75;57;51m_[38;2;77;60;49m_[38;2;77;60;50m__[38;2;77;59;49m_[38;2;76;58;48m_[38;2;75;57;47m++[38;2;77;59;49m__[38;2;78;60;50m_[38;2;79;60;50m_[38;2;79;59;50m_[38;2;80;60;51m_[38;2;78;58;49m_[38;2;75;56;48m+");
  $display("[38;2;89;88;93mjjjjjj[38;2;88;87;92mj[38;2;89;88;92mj[38;2;90;89;94mj[38;2;76;70;70m?[38;2;80;65;57m-[38;2;79;61;52m-[38;2;119;102;94mn[38;2;223;206;198ma[38;2;225;208;200mo[38;2;224;207;199maaaa[38;2;225;208;200mo[38;2;227;210;202mo[38;2;124;107;99mv[38;2;76;58;50m_[38;2;79;63;53m-[38;2;81;62;55m-[38;2;79;49;51m+[38;2;69;19;42m![38;2;79;9;46m![38;2;83;8;51mi[38;2;79;9;50mi[38;2;82;9;50mi[38;2;76;9;49m![38;2;149;111;128mY[38;2;230;212;208m*[38;2;225;208;200mo[38;2;227;210;202mo[38;2;226;209;201mo[38;2;227;208;200mo[38;2;223;208;198ma[38;2;230;206;206mo[38;2;117;75;92mr[38;2;76;10;46m![38;2;85;9;51mi[38;2;93;11;58m~[38;2;112;17;70m-[38;2;108;17;69m-[38;2;91;9;56m~[38;2;82;9;51mi[38;2;84;8;48mi[38;2;102;16;62m_[38;2;111;20;70m-[38;2;112;21;71m-[38;2;107;21;67m-[38;2;135;87;106mu[38;2;164;145;139mL[38;2;200;180;171mp[38;2;228;209;201mo[38;2;227;211;208m*[38;2;144;112;122mX[38;2;76;30;48m~[38;2;72;34;45mi[38;2;70;33;37mi[38;2;101;46;52m-[38;2;157;77;88mu[38;2;190;93;106mY[38;2;202;96;110mU[38;2;208;101;114mJ[38;2;214;111;124mL[38;2;218;119;132m0[38;2;224;124;137mO[38;2;226;125;139mO[38;2;227;127;141mZ[38;2;229;128;142mZ[38;2;230;129;143mZ[38;2;231;128;142mZZ[38;2;231;128;141mZ[38;2;229;126;140mZ[38;2;226;125;138mO[38;2;224;120;135m0[38;2;220;117;133m0[38;2;203;107;120mC[38;2;144;73;83mx[38;2;77;36;45m~[38;2;64;34;39m![38;2;66;37;40mii[38;2;64;34;40mi[38;2;184;155;162mZ[38;2;188;157;166mm[38;2;71;18;46m![38;2;81;9;53mi[38;2;82;8;52mi[38;2;79;9;50mi[38;2;85;9;53mi[38;2;97;13;62m+[38;2;99;9;62m+[38;2;110;16;70m-[38;2;111;17;70m-[38;2;95;26;57m+[38;2;83;53;53m_[38;2;79;60;51m_[38;2;79;61;50m_[38;2;81;60;52m-[38;2;81;62;51m-[38;2;80;62;52m-[38;2;80;61;53m--[38;2;80;62;52m--[38;2;80;61;52m-[38;2;79;63;52m-[38;2;67;56;52m+[38;2;62;57;61m_[38;2;61;60;64m_[38;2;61;60;65m__[38;2;60;59;64m_[38;2;59;58;63m_[38;2;60;60;67m_[38;2;61;60;69m_[38;2;61;53;61m+[38;2;71;55;55m_[38;2;80;61;54m-[38;2;81;61;52m-[38;2;81;61;53m-[38;2;80;62;52m--------[38;2;81;61;52m---[38;2;79;62;52m-[38;2;66;54;53m+[38;2;62;56;63m_[38;2;61;60;67m__[38;2;61;60;66m__[38;2;61;60;65m____[38;2;61;60;64m_[38;2;61;60;65m_[38;2;61;60;66m_[38;2;61;60;68m__[38;2;61;60;66m_[38;2;61;60;65m_[38;2;61;60;64m_[38;2;58;57;66m_[38;2;93;95;107mx[38;2;114;107;110mv[38;2;75;57;51m_[38;2;81;62;53m-[38;2;81;62;52m--[38;2;80;62;52m----[38;2;81;62;52m----[38;2;81;61;52m-[38;2;80;60;52m--[38;2;79;60;53m-");
  $display("[38;2;89;88;93mjjjjjjj[38;2;90;89;93mj[38;2;91;90;95mr[38;2;75;68;68m?[38;2;78;63;54m-[38;2;82;64;54m-[38;2;80;63;54m-[38;2;173;156;149m0[38;2;230;213;206m*[38;2;224;207;199maa[38;2;225;208;200mooo[38;2;230;213;205m*[38;2;186;169;161mm[38;2;80;63;55m-[38;2;80;61;54m-[38;2;81;61;54m-[38;2;82;60;54m-[38;2;73;41;48m~[38;2;72;14;43m![38;2;80;9;50mi[38;2;78;10;49m![38;2;80;10;49mi[38;2;76;9;47m![38;2;155;116;131mU[38;2;232;214;208m*[38;2;221;204;196ma[38;2;205;188;180md[38;2;202;185;177md[38;2;209;192;184mb[38;2;222;209;200ma[38;2;226;202;203ma[38;2;104;61;80mt[38;2;78;10;49m![38;2;83;9;51mi[38;2;82;7;51mi[38;2;101;13;64m+[38;2;105;18;69m-[38;2;89;8;55mi[38;2;83;9;51mi[38;2;84;8;49mi[38;2;98;11;61m+[38;2;112;17;73m-[38;2;112;19;72m-[38;2;109;18;68m-[38;2;114;51;80mt[38;2;147;124;123mY[38;2;169;148;140mQ[38;2;218;199;193mh[38;2;226;212;207m*[38;2;213;190;190mk[38;2;103;64;72mt[38;2;74;29;39mi[38;2;113;50;64m1[38;2;184;94;114mY[38;2;197;95;114mU[38;2;209;108;124mL[38;2;224;123;137mO[38;2;229;129;142mZ[38;2;228;130;143mZ[38;2;227;129;142mZZ[38;2;229;130;142mZ[38;2;229;128;142mZZZZZZZ[38;2;229;129;143mZ[38;2;230;129;143mZ[38;2;231;130;144mZ[38;2;233;130;145mZ[38;2;229;128;146mZ[38;2;181;103;117mU[38;2;98;47;55m-[38;2;66;34;40mi[38;2;64;36;41mi[38;2;73;47;52m+[38;2;212;186;192mb[38;2;153;112;130mY[38;2;70;8;43ml[38;2;80;8;52mi[38;2;79;9;51mi[38;2;81;9;49mi[38;2;84;9;52mi[38;2;87;11;56m~[38;2;92;12;59m~[38;2;110;16;72m-[38;2;106;18;68m-[38;2;89;35;58m_[38;2;82;59;55m-[38;2;80;60;53m---[38;2;80;60;51m_[38;2;79;59;50m_[38;2;77;57;48m_[38;2;78;58;49m_[38;2;79;59;50m_[38;2;78;58;49m__[38;2;77;61;52m_[38;2;67;55;54m+[38;2;61;56;62m+[38;2;61;61;66m_[38;2;61;60;65m_[38;2;60;59;65m_[38;2;60;59;64m_[38;2;61;59;65m_[38;2;61;60;68m_[38;2;61;59;69m_[38;2;61;53;60m+[38;2;70;56;53m+[38;2;79;62;55m-[38;2;80;61;53m-[38;2;81;61;52m-[38;2;80;62;52m----[38;2;79;62;51m-[38;2;80;62;51m-[38;2;80;62;52m--[38;2;81;61;52m--[38;2;82;62;53m-[38;2;78;61;53m-[38;2;66;54;53m+[38;2;62;56;63m_[38;2;59;58;64m___[38;2;59;58;65m_[38;2;61;60;66m_[38;2;61;60;65m___[38;2;61;60;64m_[38;2;61;60;65m_[38;2;61;60;66m_[38;2;60;59;67m_[38;2;56;55;64m+[38;2;54;53;59m+[38;2;54;53;58m+[38;2;59;58;62m+[38;2;58;57;66m_[38;2;89;92;104mr[38;2;112;107;110mu[38;2;73;58;51m_[38;2;80;62;52m-------[38;2;81;61;52m--[38;2;80;60;51m__[38;2;79;59;52m___[38;2;79;60;53m-");
  $display("[38;2;89;88;93mjjjjjj[38;2;88;87;92mj[38;2;90;89;93mj[38;2;91;89;94mj[38;2;76;68;68m?[38;2;77;62;53m-[38;2;82;64;54m-[38;2;79;61;52m-[38;2;105;88;79mj[38;2;219;201;193mh[38;2;226;209;200mo[38;2;223;206;198ma[38;2;219;202;195mh[38;2;214;198;190mk[38;2;213;196;188mk[38;2;220;203;195ma[38;2;229;212;204m*[38;2;150;133;125mU[38;2;78;60;52m_[38;2;81;61;54m-[38;2;82;61;54m-[38;2;79;59;56m-[38;2;72;30;48mi[38;2;76;11;48m![38;2;80;9;49mi[38;2;80;11;48mi[38;2;76;11;44m![38;2;162;126;137mJ[38;2;231;214;208m*[38;2;219;202;194mh[38;2;198;181;173mp[38;2;197;180;172mp[38;2;205;189;181md[38;2;223;208;200ma[38;2;221;200;200ma[38;2;103;58;77mt[38;2;79;10;49mi[38;2;83;11;53mi[38;2;79;8;50m![38;2;88;9;54mi[38;2;100;19;65m_[38;2;87;9;53mi[38;2;83;7;50mi[38;2;84;6;51mi[38;2;94;7;61m~[38;2;109;15;73m-[38;2;113;17;72m-[38;2;112;17;69m-[38;2;106;35;71m?[38;2;154;121;130mU[38;2;145;123;120mY[38;2;171;151;146m0[38;2;222;204;197ma[38;2;232;213;206m*[38;2;196;170;168mw[38;2;90;52;58m-[38;2;95;36;51m_[38;2;161;80;100mv[38;2;216;116;133mQ[38;2;233;130;146mZ[38;2;230;130;143mZ[38;2;226;130;141mZ[38;2;227;128;141mZ[38;2;227;128;142mZ[38;2;228;129;142mZ[38;2;229;129;142mZ[38;2;229;128;143mZZZ[38;2;229;128;142mZZZZZZZ[38;2;228;128;142mZ[38;2;231;128;142mZ[38;2;236;132;147mm[38;2;204;117;132mQ[38;2;94;44;56m-[38;2;63;29;41m![38;2;95;65;70m1[38;2;223;194;198mh[38;2;112;57;85mf[38;2;78;7;49m![38;2;80;9;53mi[38;2;79;9;48m![38;2;80;9;47m![38;2;81;8;48m![38;2;82;7;50mi[38;2;88;11;54m~[38;2;105;19;66m_[38;2;100;24;62m_[38;2;87;47;57m_[38;2;81;61;54m-[38;2;80;61;53m--[38;2;80;61;52m-[38;2;79;59;50m__[38;2;78;58;49m_[38;2;79;59;50m_[38;2;80;60;51m_[38;2;79;59;50m_[38;2;80;60;51m_[38;2;78;62;53m-[38;2;67;56;54m+[38;2;61;56;62m+[38;2;59;60;65m_[38;2;60;59;63m_[38;2;65;64;67m-[38;2;64;63;66m-[38;2;58;58;59m+[38;2;60;59;63m_[38;2;62;60;67m_[38;2;62;54;59m+[38;2;70;56;52m+[38;2;75;59;51m_[38;2;75;57;49m_[38;2;76;57;47m_[38;2;75;57;48m__[38;2;76;57;49m__[38;2;76;57;48m_[38;2;76;58;49m_[38;2;77;59;50m_[38;2;80;61;52m-[38;2;81;61;52m--[38;2;81;61;51m-[38;2;79;61;53m-[38;2;67;54;53m+[38;2;63;56;63m_[38;2;60;59;65m____[38;2;61;60;66m_[38;2;61;60;65m___[38;2;61;60;64m_[38;2;61;60;65m_[38;2;59;58;64m_[38;2;64;63;69m-[38;2;113;112;118mv[38;2;171;170;175mm[38;2;156;156;159m0[38;2;82;81;85mt[38;2;53;54;62m+[38;2;84;89;99mj[38;2;112;108;109mu[38;2;74;59;52m_[38;2;80;62;52m----[38;2;78;60;50m_[38;2;77;59;49m_[38;2;76;58;48m_[38;2;77;58;48m_[38;2;77;58;49m_[38;2;77;57;48m_[38;2;76;57;48m_[38;2;76;57;49m_[38;2;78;59;50m_[38;2;78;59;51m__");
  $display("[38;2;89;88;93mjjjjjjj[38;2;89;88;94mj[38;2;92;88;94mj[38;2;77;67;67m?[38;2;76;62;50m_[38;2;82;64;53m-[38;2;82;64;54m-[38;2;77;59;49m_[38;2;156;138;128mJ[38;2;232;213;203m*[38;2;212;194;186mk[38;2;183;167;159mZ[38;2;172;155;148m0[38;2;175;158;150mO[38;2;205;188;180md[38;2;229;212;204m*[38;2;224;208;199ma[38;2;123;106;98mu[38;2;75;56;49m_[38;2;79;60;53m-[38;2;79;56;56m_[38;2;73;28;49mi[38;2;73;12;47m![38;2;75;10;49m![38;2;80;10;51mi[38;2;78;16;49mi[38;2;187;153;165mZ[38;2;229;211;206m*[38;2;225;208;200mo[38;2;226;209;201mo[38;2;226;210;201mo[38;2;225;209;201mo[38;2;225;208;200mo[38;2;218;200;199mh[38;2;104;57;76mt[38;2;78;9;49m![38;2;82;10;54mi[38;2;81;8;50mi[38;2;83;7;48mi[38;2;89;12;54m~[38;2;85;10;51mi[38;2;81;8;49mi[38;2;84;8;50mi[38;2;90;7;57m~[38;2;106;14;69m_[38;2;113;16;70m-[38;2;114;18;73m-[38;2;100;23;67m_[38;2;141;95;115mc[38;2;166;142;143mL[38;2;143;124;118mY[38;2;166;147;141mQ[38;2;220;201;195mh[38;2;235;213;209m*[38;2;192;164;165mm[38;2;92;50;57m-[38;2;93;33;46m+[38;2;186;104;119mU[38;2;234;134;152mm[38;2;232;129;144mZ[38;2;228;130;142mZ[38;2;229;128;142mZZZZZZZZZZZZZZ[38;2;228;128;142mZ[38;2;228;128;143mZ[38;2;230;127;144mZ[38;2;233;134;151mm[38;2;164;93;106mz[38;2;66;21;39m![38;2;136;108;113mz[38;2;200;172;177mp[38;2;80;23;53m~[38;2;82;8;51mi[38;2;79;9;51mi[38;2;81;8;47m![38;2;79;7;48m![38;2;81;7;48m![38;2;83;5;47m![38;2;96;11;57m~[38;2;101;22;62m_[38;2;88;38;55m_[38;2;80;60;54m-[38;2;79;62;51m-[38;2;80;62;51m---[38;2;81;60;51m-[38;2;81;61;52m------[38;2;78;62;53m-[38;2;68;56;55m+[38;2;61;56;63m_[38;2;62;62;67m_[38;2;91;90;94mj[38;2;108;108;109mu[38;2;195;195;195mb[38;2;166;166;164mZ[38;2;70;69;71m?[38;2;60;58;65m_[38;2;62;55;59m+[38;2;69;55;52m+[38;2;75;60;52m_[38;2;75;59;50m_[38;2;75;57;47m+[38;2;75;56;49m__[38;2;76;57;51m__[38;2;77;57;50m_[38;2;76;56;49m_[38;2;77;57;50m_[38;2;78;58;51m_[38;2;80;60;53m-[38;2;81;61;51m-[38;2;81;61;49m_[38;2;80;61;53m-[38;2;69;54;54m+[38;2;63;56;63m_[38;2;61;59;65m_[38;2;61;60;66m____[38;2;61;60;65m_____[38;2;57;56;61m+[38;2;96;95;100mx[38;2;130;130;134mY[38;2;153;152;156mQ[38;2;158;158;161m0[38;2;124;124;128mX[38;2;55;57;63m+[38;2;81;86;95mj[38;2;112;107;107mu[38;2;75;58;50m_[38;2;80;61;51m-[38;2;80;62;51m--[38;2;79;61;51m___[38;2;80;62;51m-[38;2;80;62;52m--------");
  $display("[38;2;89;88;93mjjjjjj[38;2;88;87;92mj[38;2;89;88;93mj[38;2;92;88;95mj[38;2;77;67;68m?[38;2;76;61;51m_[38;2;81;63;52m-[38;2;82;64;54m-[38;2;80;62;52m-[38;2;91;72;63m1[38;2;203;184;175mp[38;2;229;211;203mo[38;2;221;204;197ma[38;2;215;197;190mk[38;2;222;205;197ma[38;2;225;208;200moo[38;2;227;211;203mo[38;2;212;196;188mk[38;2;106;88;80mj[38;2;76;53;50m+[38;2;73;32;48m~[38;2;76;12;45m![38;2;77;11;49m![38;2;77;13;49mi[38;2;75;11;45m![38;2;107;59;81mt[38;2;224;198;202ma[38;2;225;208;201mo[38;2;224;207;199maaa[38;2;223;207;199ma[38;2;225;208;200mo[38;2;219;201;199ma[38;2;106;58;78mt[38;2;80;9;49mi[38;2;83;11;55mi[38;2;81;8;50mi[38;2;81;7;47m![38;2;82;8;49mi[38;2;80;8;48m![38;2;79;8;48m![38;2;81;7;47m![38;2;84;6;51mi[38;2;99;12;62m+[38;2;110;17;69m-[38;2;112;16;73m-[38;2;106;18;67m_[38;2;115;56;84mf[38;2;168;140;145mQ[38;2;159;141;135mC[38;2;132;114;107mc[38;2;162;142;137mL[38;2;206;190;184mb[38;2;229;212;205m*[38;2;203;177;173mp[38;2;107;69;73mf[38;2;88;33;46m+[38;2;172;99;114mY[38;2;223;133;150mZ[38;2;226;129;144mZ[38;2;229;127;142mZ[38;2;231;127;142mZ[38;2;230;127;141mZ[38;2;230;128;140mZ[38;2;231;129;140mZ[38;2;230;129;139mZ[38;2;231;129;140mZ[38;2;232;128;142mZ[38;2;231;128;142mZ[38;2;231;128;143mZ[38;2;231;129;143mZ[38;2;230;128;143mZZ[38;2;229;128;142mZ[38;2;227;127;140mO[38;2;225;125;139mO[38;2;223;126;142mO[38;2;218;132;146mZ[38;2;194;134;145m0[38;2;84;44;57m_[38;2;187;160;166mm[38;2;145;113;124mX[38;2;70;9;41ml[38;2;83;4;48m![38;2;80;9;52mi[38;2;82;9;49mi[38;2;79;10;48m![38;2;83;8;48mi[38;2;89;8;50mi[38;2;106;19;64m_[38;2;94;31;60m_[38;2;81;56;57m-[38;2;79;62;53m-[38;2;80;62;53m-[38;2;80;62;54m--[38;2;80;62;53m-[38;2;80;61;52m-[38;2;78;58;49m_[38;2;79;57;48m_[38;2;80;57;49m_[38;2;79;58;50m_[38;2;79;60;50m_[38;2;78;61;50m_[38;2;77;61;53m_[38;2;68;56;55m+[38;2;61;56;61m+[38;2;62;62;67m_[38;2;87;86;91mj[38;2;90;90;94mj[38;2;122;122;125mz[38;2;140;140;141mJ[38;2;92;91;94mr[38;2;60;57;63m_[38;2;63;56;60m+[38;2;70;57;54m_[38;2;75;59;50m_[38;2;78;60;50m_[38;2;79;61;51m_[38;2;78;60;50m_[38;2;77;59;49m_[38;2;78;60;50m_[38;2;77;59;50m_[38;2;78;57;51m__[38;2;78;58;51m_[38;2;76;56;47m+[38;2;77;57;48m_[38;2;80;60;51m_[38;2;81;62;51m-[38;2;80;62;54m-[38;2;71;56;55m_[38;2;64;57;63m_[38;2;62;60;66m_[38;2;61;61;67m___[38;2;62;61;66m_[38;2;61;60;65m_[38;2;59;58;62m+[38;2;59;58;63m_[38;2;60;60;64m_[38;2;61;60;64m_[38;2;61;60;65m_[38;2;65;64;69m-[38;2;72;71;77m?[38;2;75;74;79m1[38;2;72;71;76m?[38;2;69;68;72m?[38;2;59;58;65m_[38;2;82;82;91mf[38;2;114;104;106mu[38;2;75;58;51m_[38;2;80;62;52m-[38;2;81;62;53m-[38;2;81;63;53m-[38;2;80;63;53m-[38;2;81;63;53m-[38;2;81;62;52m-[38;2;79;60;50m_[38;2;78;60;48m_[38;2;80;61;51m-[38;2;81;61;53m-[38;2;81;62;52m-[38;2;80;62;52m---[38;2;79;61;51m_");
  $display("[38;2;89;88;93mjjjjjjj[38;2;90;89;94mj[38;2;93;89;96mr[38;2;77;66;69m?[38;2;75;59;53m_[38;2;79;61;51m_[38;2;81;63;53m-[38;2;82;64;54m-[38;2;76;58;49m_[38;2;133;114;107mc[38;2;228;209;202mo[38;2;226;207;200moo[38;2;225;208;200mo[38;2;224;207;199maa[38;2;224;208;201mo[38;2;228;215;205m*[38;2;194;178;169mq[38;2;82;54;58m-[38;2;72;15;44m![38;2;85;11;52mi[38;2;77;12;50mi[38;2;79;12;48mi[38;2;73;14;43m![38;2;165;127;139mC[38;2;234;212;210m*[38;2;224;207;199maaaa[38;2;223;207;199ma[38;2;225;208;200mo[38;2;223;205;203ma[38;2;112;65;84mj[38;2;80;9;49mi[38;2;82;11;55mi[38;2;81;9;50mi[38;2;79;8;47m![38;2;79;8;48m![38;2;78;7;47m![38;2;79;8;48m![38;2;81;7;48m![38;2;81;7;49m![38;2;89;9;54mi[38;2;106;17;67m_[38;2;113;18;72m-[38;2;114;18;72m-[38;2;101;28;66m-[38;2;150;110;126mY[38;2;166;147;146mQ[38;2;150;131;124mU[38;2;147;128;122mY[38;2;156;139;133mC[38;2;169;150;144mQ[38;2;204;183;178md[38;2;216;193;189mk[38;2;143;117;117mX[38;2;87;43;51m_[38;2;127;74;85mr[38;2;195;145;155mZ[38;2;207;154;163mw[38;2;208;146;156mm[38;2;211;143;153mZ[38;2;210;140;149mZ[38;2;209;139;147mZ[38;2;210;135;145mO[38;2;210;132;143mO[38;2;213;133;146mO[38;2;214;134;149mZ[38;2;214;136;150mZ[38;2;213;138;151mZ[38;2;209;139;151mZ[38;2;206;141;152mZ[38;2;211;151;160mw[38;2;211;160;167mq[38;2;215;176;181md[38;2;198;169;173mq[38;2;237;221;223mM[38;2;182;167;172mm[38;2;106;74;82mj[38;2;195;160;171mw[38;2;81;32;55m+[38;2;86;28;60m+[38;2;111;76;105mx[38;2;116;99;122mv[38;2;116;96;121mv[38;2;113;96;122mv[38;2;115;95;122mv[38;2;117;95;123mv[38;2;121;97;126mv[38;2;117;100;127mv[38;2;114;106;125mc[38;2;115;105;122mvv[38;2;115;105;123mvv[38;2;116;105;122mv[38;2;117;105;121mv[38;2;112;99;109mu[38;2;101;86;91mr[38;2;90;72;73mt[38;2;79;60;54m-[38;2;74;55;44m+[38;2;75;56;47m+[38;2;76;60;53m_[38;2;67;56;53m+[38;2;60;56;58m+[38;2;70;69;78m?[38;2;106;101;113mu[38;2;121;115;130mz[38;2;115;106;129mc[38;2;119;110;133mz[38;2;115;106;127mc[38;2;115;104;125mv[38;2;117;105;124mc[38;2;116;106;117mv[38;2;103;91;94mx[38;2;81;64;58m-[38;2;79;61;49m_[38;2;78;60;50m_[38;2;77;59;49m__[38;2;77;59;50m_[38;2;76;58;51m_[38;2;74;57;47m+[38;2;77;59;51m_[38;2;86;71;68m1[38;2;102;90;94mr[38;2;116;103;116mv[38;2;119;106;121mc[38;2;119;105;124mc[38;2;117;104;123mv[38;2;116;104;124mv[38;2;116;105;126mc[38;2;116;105;125mccc[38;2;116;106;127mc[38;2;113;107;126mc[38;2;102;98;111mn[38;2;83;81;89mf[38;2;65;64;70m-[38;2;58;57;63m+[38;2;60;59;64m_[38;2;59;58;62m+[38;2;59;57;61m+[38;2;72;69;76m?[38;2;89;86;97mj[38;2;105;100;114mu[38;2;116;106;123mc[38;2;118;110;129mz[38;2;126;114;133mX[38;2;120;104;123mc[38;2;120;105;123mc[38;2;121;105;124mcc[38;2;122;105;124mc[38;2;122;106;123mc[38;2;120;107;120mc[38;2;112;101;109mu[38;2;99;85;87mj[38;2;83;68;58m?[38;2;76;58;46m_[38;2;77;58;49m_[38;2;78;60;50m__[38;2;77;59;50m_[38;2;77;59;49m_");
  $display("[38;2;89;88;93mjjjjjjj[38;2;90;89;94mj[38;2;93;89;96mr[38;2;79;69;71m?[38;2;70;54;48m+[38;2;75;56;47m+[38;2;77;59;49m_[38;2;78;60;51m_[38;2;77;59;50m_[38;2;81;62;55m-[38;2;192;173;166mw[38;2;228;211;203mo[38;2;224;206;199ma[38;2;224;207;199maaa[38;2;224;207;200ma[38;2;224;209;200mo[38;2;230;214;205m*[38;2;174;149;150m0[38;2;76;23;48mi[38;2;85;10;51mi[38;2;84;11;52mi[38;2;80;10;46m![38;2;96;41;64m-[38;2;217;188;192mk[38;2;228;210;202mo[38;2;224;207;198ma[38;2;224;207;199maaa[38;2;223;207;198ma[38;2;225;208;200mo[38;2;224;205;205mo[38;2;115;68;88mj[38;2;77;10;49m![38;2;81;11;54mi[38;2;82;8;50mi[38;2;81;8;48m![38;2;79;8;48m!![38;2;78;7;47m![38;2;79;8;48m![38;2;79;8;49m![38;2;83;7;50mi[38;2;95;12;59m+[38;2;109;20;71m-[38;2;117;18;74m?[38;2;106;20;68m-[38;2;119;63;91mj[38;2;170;142;147mQ[38;2;154;134;129mJ[38;2;135;117;107mz[38;2;155;135;129mJ[38;2;162;143;137mL[38;2;157;139;132mC[38;2;168;151;144mQ[38;2;196;178;173mq[38;2;186;162;162mm[38;2;119;89;95mn[38;2;94;62;72m1[38;2;127;98;108mv[38;2;196;177;184mp[38;2;240;232;234m&[38;2;244;239;241m8[38;2;239;234;236m&[38;2;230;226;227mM[38;2;193;187;187md[38;2;230;223;223mM[38;2;232;227;227mM[38;2;234;229;230mW[38;2;236;233;233m&[38;2;227;222;224mM[38;2;209;206;207ma[38;2;246;247;247mB[38;2;247;252;250m@[38;2;255;255;255m$[38;2;216;212;214mo[38;2;170;152;159mO[38;2;76;50;57m_[38;2;165;131;141mC[38;2;127;79;101mn[38;2;74;10;45m![38;2;119;95;117mv[38;2;128;129;144mU[38;2;127;123;130mX[38;2;160;159;119mC[38;2;168;166;117mL[38;2;167;165;117mL[38;2;165;166;116mL[38;2;164;165;116mL[38;2;164;165;117mL[38;2;162;165;116mL[38;2;162;164;117mL[38;2;160;165;117mL[38;2;159;165;117mL[38;2;157;164;116mCC[38;2;147;149;119mJ[38;2;132;129;128mY[38;2;126;119;137mX[38;2;125;117;141mX[38;2;121;113;123mz[38;2;101;90;90mr[38;2;80;64;56m-[38;2;76;60;51m_[38;2;66;54;48m+[38;2;69;62;69m-[38;2;117;115;128mz[38;2;129;124;140mY[38;2;125;124;130mX[38;2;143;162;115mJ[38;2;144;163;117mJ[38;2;142;165;113mJ[38;2;144;165;118mC[38;2;139;152;121mU[38;2;124;120;134mX[38;2;131;125;141mY[38;2;108;100;108mn[38;2;79;60;51m_[38;2;81;61;50m-[38;2;81;62;52m-[38;2;80;61;52m-[38;2;79;61;52m-[38;2;77;60;51m_[38;2;92;78;74mt[38;2;116;107;116mv[38;2;129;118;139mY[38;2;127;119;138mY[38;2;122;129;129mX[38;2;126;154;119mU[38;2;128;165;114mU[38;2;127;165;115mU[38;2;125;165;115mU[38;2;124;165;115mU[38;2;124;165;114mU[38;2;123;165;114mUU[38;2;122;163;116mU[38;2;122;139;125mY[38;2;127;121;137mY[38;2;129;120;139mY[38;2;120;114;131mz[38;2;92;90;100mr[38;2;65;61;71m-[38;2;74;71;78m1[38;2;108;101;115mu[38;2;127;118;136mX[38;2;130;118;140mY[38;2;123;125;130mX[38;2;115;148;120mX[38;2;108;165;113mY[38;2;106;164;114mY[38;2;107;165;116mY[38;2;108;164;117mY[38;2;108;163;116mY[38;2;106;164;115mY[38;2;104;164;116mY[38;2;105;163;117mY[38;2;110;144;122mX[38;2;123;122;133mX[38;2;131;119;140mY[38;2;127;115;132mX[38;2;106;95;99mx[38;2;82;65;60m?[38;2;76;58;47m_[38;2;79;60;49m_[38;2;78;60;50m__");
  $display("[38;2;89;88;93mjjjjjjj[38;2;90;89;94mj[38;2;93;89;96mr[38;2;79;69;72m?[38;2;74;58;52m_[38;2;79;61;53m-[38;2;80;61;54m-[38;2;78;59;52m_[38;2;80;61;54m-[38;2;77;58;51m_[38;2;133;116;108mz[38;2;226;212;203mo[38;2;224;209;200mo[38;2;224;207;199maaaa[38;2;225;208;200moo[38;2;230;212;205m*[38;2;140;100;113mc[38;2;75;11;42m![38;2;82;10;48mi[38;2;68;5;38ml[38;2;123;78;96mx[38;2;232;209;208m*[38;2;225;208;200mo[38;2;224;207;199maaaa[38;2;223;208;197ma[38;2;225;208;199ma[38;2;224;206;206mo[38;2;117;71;92mr[38;2;77;10;49m![38;2;80;11;51mi[38;2;80;9;49mi[38;2;81;9;49mi[38;2;80;9;49mii[38;2;78;7;47m![38;2;79;8;48m![38;2;80;8;48m![38;2;79;8;47m![38;2;80;8;48m![38;2;99;17;63m+[38;2;114;19;69m-[38;2;112;20;69m-[38;2;100;27;65m-[38;2;149;106;120mX[38;2;166;145;142mQ[38;2;142;121;112mX[38;2;137;116;108mz[38;2;157;138;131mC[38;2;165;146;139mL[38;2;161;143;136mC[38;2;157;138;131mC[38;2;166;146;140mL[38;2;189;168;165mw[38;2;176;152;151m0[38;2;131;101;105mv[38;2;94;59;69m1[38;2;110;80;92mr[38;2;158;137;149mL[38;2;199;185;195mb[38;2;221;215;219m*[38;2;207;204;204mh[38;2;253;252;253m$[38;2;252;251;251m@[38;2;251;251;251m@[38;2;252;252;252m$[38;2;241;240;243m8[38;2;205;196;202mk[38;2;233;222;229mM[38;2;214;204;209ma[38;2;180;163;169mm[38;2;113;80;91mr[38;2;71;29;42mi[38;2;147;110;118mX[38;2;182;153;160mZ[38;2;75;18;46mi[38;2;86;16;56m~[38;2;125;106;126mz[38;2;126;121;140mY[38;2;115;114;103mv[38;2;232;232;78mq[38;2;254;255;71mb[38;2;248;254;70md[38;2;244;255;69md[38;2;244;255;68md[38;2;245;255;68md[38;2;242;255;68md[38;2;238;255;69mp[38;2;236;255;69mp[38;2;232;255;69mp[38;2;228;255;70mp[38;2;223;255;69mq[38;2;216;251;70mq[38;2;204;235;73mm[38;2;181;205;88m0[38;2;146;154;105mU[38;2;124;118;129mz[38;2;129;122;144mY[38;2;120;111;124mc[38;2;87;75;68m1[38;2;65;53;47m+[38;2;106;96;110mn[38;2;131;124;143mY[38;2;118;112;125mc[38;2;145;177;91mU[38;2;185;255;67mZ[38;2;180;255;69mZ[38;2;177;255;64mZ[38;2;174;255;71mZ[38;2;169;245;70mO[38;2;120;140;99mz[38;2;126;114;139mX[38;2;129;124;136mY[38;2;98;83;83mj[38;2;78;59;46m_[38;2;80;62;51m-[38;2;80;61;53m-[38;2;79;60;52m_[38;2;102;90;93mr[38;2;129;121;138mY[38;2;129;119;137mY[38;2;118;133;119mz[38;2;125;191;92mU[38;2;127;234;72mC[38;2;128;252;67mL[38;2;127;255;66mL[38;2;126;255;66mL[38;2;122;255;65mL[38;2;119;255;64mC[38;2;117;255;65mC[38;2;112;255;64mC[38;2;109;255;66mC[38;2;107;254;69mC[38;2;103;244;70mJ[38;2;101;215;78mY[38;2;109;155;105mz[38;2;123;117;134mX[38;2;131;122;142mY[38;2;115;113;122mc[38;2;125;116;132mX[38;2;130;121;141mY[38;2;117;125;120mz[38;2;95;180;91mz[38;2;80;228;76mY[38;2;73;251;66mY[38;2;67;255;62mY[38;2;67;255;65mY[38;2;63;255;64mX[38;2;59;255;61mX[38;2;57;255;61mX[38;2;54;255;66mX[38;2;52;255;65mX[38;2;47;255;63mz[38;2;51;247;69mz[38;2;59;223;73mc[38;2;81;169;96mc[38;2;118;120;131mz[38;2;132;122;140mY[38;2;122;115;126mz[38;2;90;74;72mt[38;2;79;60;48m_[38;2;80;62;51m-[38;2;80;61;52m-");
  $display("[38;2;89;88;93mjjjjjjjj[38;2;91;88;93mj[38;2;77;67;68m?[38;2;75;59;53m_[38;2;79;61;53m-[38;2;77;59;52m_[38;2;75;56;49m_[38;2;76;57;50m_[38;2;79;61;53m-[38;2;82;65;57m-[38;2;188;173;164mw[38;2;227;212;203mo[38;2;224;207;199maaaaaa[38;2;229;211;203mo[38;2;211;183;186mb[38;2;106;67;81mf[38;2;116;67;88mj[38;2;139;93;110mv[38;2;188;158;162mZ[38;2;229;212;206m*[38;2;225;209;201mo[38;2;225;207;200ma[38;2;222;205;197ma[38;2;221;204;196ma[38;2;222;205;197ma[38;2;224;208;198ma[38;2;226;209;201mo[38;2;226;207;207mo[38;2;119;73;94mr[38;2;77;10;48m![38;2;80;10;51mi[38;2;78;8;49m![38;2;80;9;49miii[38;2;79;8;48m!![38;2;80;8;48m!![38;2;80;7;48m![38;2;91;10;55m~[38;2;109;19;67m-[38;2;112;18;69m-[38;2;108;17;67m-[38;2;113;47;79mt[38;2;167;135;136mC[38;2;163;144;136mL[38;2;141;122;114mX[38;2;140;121;112mX[38;2;162;143;134mC[38;2;164;145;136mL[38;2;164;144;135mL[38;2;161;143;134mC[38;2;156;139;131mC[38;2;162;146;139mL[38;2;185;168;162mm[38;2;196;175;172mq[38;2;172;145;147mQ[38;2;131;98;104mv[38;2;104;65;75mt[38;2;98;58;70m1[38;2;107;72;82mj[38;2;129;98;107mv[38;2;140;109;118mz[38;2;141;110;120mz[38;2;135;105;114mc[38;2;119;85;99mn[38;2;99;55;71m1[38;2;95;47;64m-[38;2;85;41;56m_[38;2;87;43;56m_[38;2;110;67;76mf[38;2;171;143;144mQ[38;2;236;209;212m*[38;2;118;78;91mr[38;2;77;8;41m![38;2;86;18;56m~[38;2;123;106;125mc[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;230;78mq[38;2;251;255;71mb[38;2;245;252;70md[38;2;243;254;70md[38;2;231;242;71mq[38;2;189;197;67mQ[38;2;186;197;71mQ[38;2;185;198;72mQ[38;2;183;197;71mL[38;2;181;198;70mL[38;2;187;210;67mQ[38;2;209;239;68mm[38;2;221;255;69mq[38;2;216;254;70mq[38;2;215;255;65mw[38;2;211;253;69mw[38;2;172;199;85mQ[38;2;121;120;116mz[38;2;129;122;137mY[38;2;123;114;127mz[38;2;99;91;97mr[38;2;129;121;137mY[38;2;124;116;135mX[38;2;124;139;98mz[38;2;182;247;72mZ[38;2;182;254;65mZ[38;2;176;253;69mZ[38;2;177;253;68mZ[38;2;173;253;65mO[38;2;171;255;65mO[38;2;156;219;78mQ[38;2;112;119;111mv[38;2;128;121;140mY[38;2;123;115;132mz[38;2;82;69;59m?[38;2;75;59;47m_[38;2;75;59;49m_[38;2;94;80;80mf[38;2;127;123;136mY[38;2;128;116;140mY[38;2;114;141;99mc[38;2;134;236;74mL[38;2;136;255;64mQ[38;2;131;255;65mL[38;2;129;254;67mL[38;2;123;243;67mC[38;2;105;198;67mz[38;2;97;168;68mv[38;2;94;153;73mu[38;2;92;158;73mu[38;2;92;183;66mv[38;2;102;223;69mY[38;2;106;255;63mJ[38;2;104;253;65mJ[38;2;100;255;65mJ[38;2;100;252;68mJ[38;2;98;186;84mz[38;2;119;116;126mz[38;2;130;123;140mY[38;2;128;120;139mY[38;2;105;127;112mv[38;2;85;220;76mX[38;2;76;255;61mY[38;2;74;255;64mY[38;2;72;254;66mY[38;2;72;249;66mY[38;2;68;204;66mv[38;2;67;171;70mn[38;2;68;154;73mx[38;2;66;155;73mx[38;2;60;176;69mn[38;2;55;214;65mv[38;2;50;253;63mz[38;2;46;255;65mz[38;2;45;255;64mz[38;2;40;255;63mz[38;2;57;204;81mv[38;2;112;119;119mc[38;2;128;123;143mY[38;2;124;113;125mz[38;2;84;68;61m?[38;2;80;60;51m_[38;2;81;61;54m-");
  $display("[38;2;89;88;93mjjjjjjj[38;2;88;89;93mj[38;2;90;89;89mj[38;2;77;69;64m?[38;2;74;61;52m_[38;2;73;57;48m+[38;2;82;65;57m-[38;2;95;78;70mt[38;2;94;77;69mt[38;2;88;71;63m1[38;2;79;62;54m-[38;2;110;93;85mx[38;2;216;199;191mh[38;2;225;208;200mo[38;2;224;207;199maa[38;2;224;208;199ma[38;2;226;209;201mo[38;2;224;207;199ma[38;2;225;208;200mo[38;2;204;188;183md[38;2;196;179;175mp[38;2;188;170;166mw[38;2;209;190;186mb[38;2;212;194;187mk[38;2;210;191;185mb[38;2;216;197;191mk[38;2;224;207;199ma[38;2;215;198;190mk[38;2;197;180;172mp[38;2;203;186;178md[38;2;224;206;199ma[38;2;227;209;202mo[38;2;228;210;208m*[38;2;118;74;93mr[38;2;75;9;46m![38;2;83;10;51mi[38;2;81;8;51mi[38;2;80;9;51mi[38;2;80;9;49mii[38;2;79;8;48m![38;2;80;8;48m!!![38;2;80;9;48m![38;2;81;7;49m![38;2;98;14;61m+[38;2;110;19;71m-[38;2;113;18;73m-[38;2;106;19;68m-[38;2;132;80;101mn[38;2;166;145;144mQ[38;2;155;139;132mC[38;2;138;119;112mz[38;2;157;138;132mC[38;2;164;145;138mL[38;2;164;144;137mLL[38;2;163;143;136mLL[38;2;158;139;132mC[38;2;159;141;133mC[38;2;178;160;152mO[38;2;208;188;182mb[38;2;221;198;194mh[38;2;208;181;180md[38;2;184;154;157mZ[38;2;164;132;137mC[38;2;156;123;128mU[38;2;157;124;129mU[38;2;155;124;129mU[38;2;158;128;135mJ[38;2;170;138;145mQ[38;2;179;148;153mO[38;2;189;160;163mm[38;2;202;173;176mp[38;2;208;175;182md[38;2;197;161;172mw[38;2;141;97;115mc[38;2;79;20;47mi[38;2;83;10;47mi[38;2;83;17;55m~[38;2;123;106;125mc[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;229;78mq[38;2;251;254;70md[38;2;245;251;70md[38;2;245;255;71md[38;2;208;219;75mZ[38;2;100;94;99mx[38;2;110;105;123mv[38;2;112;106;123mv[38;2;115;108;124mc[38;2;114;107;123mv[38;2;110;103;117mv[38;2;110;109;92mn[38;2;164;186;68mJ[38;2;217;252;74mq[38;2;211;252;69mw[38;2;208;253;67mw[38;2;212;255;70mq[38;2;161;186;84mC[38;2;115;112;127mc[38;2;129;121;139mY[38;2;130;123;137mY[38;2;126;120;141mY[38;2;114;118;115mc[38;2;171;220;79m0[38;2;186;255;70mm[38;2;179;254;65mZ[38;2;180;252;69mZ[38;2;172;248;69mO[38;2;172;254;67mO[38;2;169;252;71mO[38;2;170;255;70mZ[38;2;138;180;87mU[38;2;115;112;127mc[38;2;130;125;141mY[38;2;109;102;107mu[38;2;73;58;47m+[38;2;73;57;47m+[38;2;111;101;108mu[38;2;129;124;140mY[38;2;116;108;123mc[38;2;122;200;82mU[38;2;140;255;65mQ[38;2;134;253;70mQ[38;2;131;254;67mL[38;2;130;247;72mL[38;2;94;134;79mn[38;2;107;99;114mu[38;2;117;109;136mz[38;2;122;109;133mz[38;2;120;110;133mz[38;2;116;105;127mc[38;2;92;103;96mx[38;2;96;199;70mz[38;2;104;255;66mJ[38;2;101;255;64mJ[38;2;98;255;62mJ[38;2;97;254;67mJ[38;2;98;142;94mv[38;2;129;115;138mX[38;2;120;112;127mz[38;2;90;169;84mv[38;2;79;255;62mY[38;2;78;252;68mY[38;2;76;253;67mY[38;2;74;253;65mY[38;2;72;158;72mx[38;2;103;97;112mn[38;2;121;108;129mz[38;2;125;110;133mz[38;2;124;110;133mz[38;2;119;106;128mc[38;2;98;100;103mx[38;2;60;173;69mx[38;2;47;255;62mz[38;2;44;255;62mz[38;2;41;255;63mz[38;2;34;255;65mc[38;2;67;167;84mu[38;2;122;112;134mz[38;2;131;123;141mY[38;2;103;91;91mr[38;2;79;63;48m_[38;2;84;64;55m-");
  $display("[38;2;89;88;93mjjjjjjj[38;2;88;89;93mj[38;2;91;89;90mj[38;2;77;68;64m?[38;2;80;66;58m-[38;2;149;132;124mU[38;2;199;181;173mp[38;2;216;199;191mh[38;2;212;195;187mk[38;2;203;186;178md[38;2;195;178;170mq[38;2;166;149;141mQ[38;2;200;183;175mp[38;2;227;210;202mo[38;2;226;209;201mo[38;2;225;208;200mo[38;2;224;207;199ma[38;2;216;198;190mk[38;2;226;208;200mo[38;2;217;200;192mh[38;2;172;154;148m0[38;2;210;193;186mb[38;2;193;178;170mq[38;2;210;195;187mk[38;2;225;206;200ma[38;2;221;202;195ma[38;2;215;195;189mk[38;2;208;190;183mb[38;2;205;188;180md[38;2;203;186;178md[38;2;211;194;186mk[38;2;213;196;188mk[38;2;217;199;192mh[38;2;223;203;203ma[38;2;136;96;111mv[38;2;73;20;48mi[38;2;80;17;50mi[38;2;77;10;47m![38;2;74;6;44ml[38;2;75;5;44ml[38;2;79;8;48m![38;2;80;9;49mi[38;2;80;8;48m!![38;2;79;7;47m![38;2;79;8;48m![38;2;79;8;49m![38;2;88;8;54mi[38;2;105;18;67m_[38;2;112;20;72m-[38;2;112;19;72m-[38;2;99;29;67m-[38;2;144;108;122mX[38;2;164;146;143mQ[38;2;136;120;114mz[38;2;137;120;114mz[38;2;157;141;135mC[38;2;163;144;137mL[38;2;163;143;136mLLL[38;2;162;143;136mLL[38;2;161;142;134mC[38;2;157;139;131mC[38;2;168;149;142mQ[38;2;190;171;165mw[38;2;200;181;176mp[38;2;203;183;180md[38;2;202;182;179mp[38;2;200;180;177mp[38;2;199;180;176mp[38;2;191;172;169mw[38;2;176;159;156mO[38;2;145;120;123mY[38;2;110;67;86mj[38;2;100;43;75m?[38;2;89;26;61m+[38;2;81;11;49mi[38;2;79;6;45m![38;2;82;9;49mi[38;2;80;7;48m![38;2;80;13;53mi[38;2;123;106;125mc[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;229;78mq[38;2;251;254;70md[38;2;245;251;70md[38;2;245;255;71md[38;2;209;220;76mZ[38;2;115;108;113mv[38;2;128;123;141mY[38;2;122;116;131mz[38;2;96;90;103mx[38;2;103;98;108mn[38;2;127;120;138mY[38;2;124;117;136mX[38;2;107;104;100mn[38;2;203;232;73mZ[38;2;213;254;71mq[38;2;208;252;72mw[38;2;207;255;68mw[38;2;188;230;73mO[38;2;113;115;112mv[38;2;126;121;135mX[38;2;131;120;142mY[38;2;116;112;126mc[38;2;148;181;82mU[38;2;192;255;71mm[38;2;183;253;67mZ[38;2;182;255;70mZ[38;2;161;218;71mL[38;2;99;134;59mx[38;2;173;248;69mO[38;2;168;253;70mO[38;2;167;254;65mO[38;2;164;247;72mO[38;2;119;145;95mz[38;2;123;114;137mX[38;2;129;124;139mY[38;2;96;86;84mj[38;2;72;58;53m_[38;2;113;101;108mu[38;2;130;124;142mY[38;2;113;106;117mv[38;2;119;193;73mY[38;2;140;255;68mQ[38;2;135;252;70mQ[38;2;131;254;66mL[38;2;127;249;68mL[38;2;109;160;87mc[38;2;124;118;127mz[38;2;127;116;138mX[38;2;127;118;138mX[38;2;127;120;140mY[38;2;131;120;141mY[38;2;123;115;136mX[38;2;102;120;104mu[38;2;93;146;83mu[38;2;90;143;83mn[38;2;88;145;82mn[38;2;91;147;84mu[38;2;102;122;104mu[38;2;125;117;136mX[38;2;118;109;127mc[38;2;85;162;79mu[38;2;81;255;64mU[38;2;78;253;66mY[38;2;73;254;64mY[38;2;73;254;67mY[38;2;77;181;79mv[38;2;116;119;125mz[38;2;128;116;137mX[38;2;130;117;141mY[38;2;129;118;141mY[38;2;130;121;142mY[38;2;131;116;141mY[38;2;98;116;109mu[38;2;74;145;85mn[38;2;69;144;79mx[38;2;68;144;83mx[38;2;69;146;80mx[38;2;85;132;104mu[38;2;126;119;133mX[38;2;135;128;145mU[38;2;80;72;78m1[38;2;39;31;28mI[38;2;40;30;30mI");
  $display("[38;2;90;89;94mjjjjjjj[38;2;90;90;94mj[38;2;93;90;92mj[38;2;74;65;61m-[38;2;123;108;100mv[38;2;231;214;205m*[38;2;228;211;203mo[38;2;226;209;201moo[38;2;227;210;202mo[38;2;228;211;203mo[38;2;229;212;204m*[38;2;225;208;200mo[38;2;200;183;175mp[38;2;210;193;185mb[38;2;220;203;195ma[38;2;203;185;178md[38;2;212;193;187mk[38;2;223;204;197ma[38;2;186;167;161mm[38;2;141;123;116mX[38;2;163;146;138mL[38;2;176;159;151mO[38;2;192;174;166mw[38;2;212;193;186mk[38;2;213;194;187mk[38;2;215;196;189mk[38;2;220;202;194mh[38;2;225;208;200mo[38;2;221;204;196ma[38;2;217;200;192mh[38;2;213;198;188mk[38;2;217;199;192mh[38;2;221;200;197ma[38;2;211;188;188mb[38;2;196;173;173mq[38;2;192;165;169mw[38;2;179;148;157mO[38;2;157;121;133mU[38;2;125;81;98mn[38;2;81;24;53m~[38;2;78;7;47m![38;2;81;8;49mi[38;2;80;8;48m!!![38;2;81;7;50mi[38;2;80;6;50m![38;2;92;11;57m~[38;2;109;19;68m-[38;2;116;18;72m-[38;2;111;18;69m-[38;2;107;41;75m1[38;2;161;127;136mJ[38;2;159;146;139mL[38;2;138;120;112mz[38;2;138;123;115mX[38;2;158;139;132mC[38;2;163;143;136mLLL[38;2;163;144;137mLLL[38;2;164;144;137mL[38;2;163;143;136mL[38;2;161;141;134mC[38;2;160;140;133mC[38;2;158;139;134mC[38;2;159;140;135mC[38;2;158;139;134mC[38;2;152;133;127mU[38;2;138;118;114mz[38;2;151;134;127mU[38;2;131;104;103mv[38;2;75;13;47m![38;2;80;9;51mi[38;2;80;8;50mi[38;2;82;8;50mi[38;2;81;9;50mi[38;2;80;9;49mi[38;2;79;7;47m![38;2;79;14;52mi[38;2;123;106;125mc[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;230;78mq[38;2;251;255;71mb[38;2;245;251;70md[38;2;245;255;71md[38;2;208;218;77mZ[38;2;110;103;112mu[38;2;123;118;140mX[38;2;122;114;138mX[38;2;112;105;123mv[38;2;114;106;127mc[38;2;123;116;137mX[38;2;120;112;136mz[38;2;129;134;95mz[38;2;210;242;73mw[38;2;212;253;69mw[38;2;208;252;70mw[38;2;210;255;70mw[38;2;182;220;72m0[38;2;109;110;112mv[38;2;127;122;138mY[38;2;123;114;136mX[38;2;128;143;101mX[38;2;190;248;71mZ[38;2;189;253;69mm[38;2;184;253;66mZ[38;2;181;252;69mZ[38;2;119;142;83mv[38;2;96;91;105mx[38;2;138;186;76mU[38;2;174;255;68mZ[38;2;168;252;68mO[38;2;165;255;69mO[38;2;151;224;74mL[38;2;112;120;112mv[38;2;128;118;142mY[38;2;125;117;130mX[38;2;90;83;87mf[38;2;101;92;99mx[38;2;129;124;135mY[38;2;126;114;137mX[38;2;100;120;89mn[38;2;126;221;71mJ[38;2;138;255;68mQ[38;2;131;255;66mL[38;2;129;253;68mL[38;2;127;252;71mL[38;2;119;226;76mJ[38;2;116;191;89mY[38;2;117;165;104mY[38;2;119;143;114mX[38;2;120;128;126mX[38;2;124;119;129mX[38;2;126;112;138mX[38;2;125;110;138mX[38;2;124;113;139mX[38;2;127;113;139mX[38;2;126;113;137mX[38;2;136;126;144mU[38;2;132;125;139mY[38;2;125;117;135mX[38;2;95;112;101mn[38;2;78;203;67mc[38;2;81;255;67mU[38;2;76;255;65mY[38;2;72;254;64mY[38;2;69;255;67mY[38;2;76;230;76mX[38;2;82;197;85mz[38;2;91;172;99mz[38;2;105;147;114mz[38;2;115;130;123mz[38;2;123;120;132mX[38;2;127;115;137mX[38;2;130;109;138mX[38;2;130;112;138mX[38;2;129;114;137mX[38;2;128;114;136mX[38;2;122;110;129mz[38;2;103;99;110mn[38;2;63;62;68m-[38;2;6;6;7m.[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;94;92;95mr[38;2;94;91;95mr[38;2;93;91;94mr[38;2;93;90;94mr[38;2;92;90;93mj[38;2;92;90;94mr[38;2;91;90;93mj[38;2;88;88;91mj[38;2;88;86;86mf[38;2;72;62;57m_[38;2;173;158;150mO[38;2;228;211;203mo[38;2;224;207;199maaaaaa[38;2;225;208;200mo[38;2;215;198;190mk[38;2;167;150;142mQ[38;2;168;151;143mQ[38;2;179;160;154mO[38;2;186;167;162mm[38;2;174;155;150m0[38;2;163;144;139mL[38;2;152;132;125mU[38;2;148;129;122mU[38;2;161;141;134mC[38;2;169;150;143mQ[38;2;199;180;173mp[38;2;221;202;195ma[38;2;223;203;196ma[38;2;222;204;197ma[38;2;228;211;203moo[38;2;226;209;201mo[38;2;222;204;196ma[38;2;216;198;191mk[38;2;210;193;185mb[38;2;214;198;189mk[38;2;226;211;202mo[38;2;228;212;204mo[38;2;228;213;204m*[38;2;232;215;207m*[38;2;232;214;210m*[38;2;185;154;164mZ[38;2;88;31;59m+[38;2;80;9;47m![38;2;82;9;50mi[38;2;81;8;49mi[38;2;80;8;47m![38;2;82;7;50mi[38;2;79;8;50m![38;2;82;8;51mi[38;2;94;14;59m+[38;2;111;18;69m-[38;2;117;17;72m-[38;2;105;19;67m_[38;2;113;57;85mf[38;2;163;138;140mL[38;2;160;141;132mC[38;2;151;130;124mU[38;2;170;150;144mQ[38;2;163;143;136mL[38;2;162;142;135mC[38;2;163;143;136mL[38;2;163;144;137mLLL[38;2;164;144;137mL[38;2;163;143;136mLLL[38;2;163;144;137mL[38;2;155;136;129mJ[38;2;146;127;120mY[38;2;140;121;114mX[38;2;143;124;116mX[38;2;166;149;139mQ[38;2;149;122;120mY[38;2;81;24;52m~[38;2;79;12;49mi[38;2;79;10;47m![38;2;79;10;48m![38;2;80;10;49mi[38;2;79;8;49m![38;2;79;7;48m![38;2;80;14;52mi[38;2;123;106;125mc[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;230;78mq[38;2;251;255;71mb[38;2;245;251;70md[38;2;244;254;71md[38;2;218;229;73mm[38;2;147;148;96mY[38;2;153;157;109mJ[38;2;155;157;111mJ[38;2;154;158;107mJ[38;2;153;157;112mJ[38;2;157;164;103mJ[38;2;174;188;92mQ[38;2;207;238;72mm[38;2;215;253;72mq[38;2;211;253;69mw[38;2;212;255;70mq[38;2;205;246;70mm[38;2;128;141;85mc[38;2;115;111;128mc[38;2;128;118;140mY[38;2;116;120;109mc[38;2;178;223;77m0[38;2;190;255;69mm[38;2;186;252;68mZ[38;2;187;255;70mm[38;2;149;197;70mJ[38;2;105;103;112mu[38;2;127;115;141mX[38;2;103;116;92mn[38;2;161;232;70mQ[38;2;167;255;66mO[38;2;166;252;69mO[38;2;162;255;70mO[38;2;135;187;84mU[38;2;116;111;124mc[38;2;131;121;139mY[38;2;117;113;126mc[38;2;90;89;95mj[38;2;109;105;111mu[38;2;129;120;137mY[38;2;121;114;132mz[38;2;99;111;99mn[38;2;108;167;70mc[38;2;121;226;66mU[38;2;126;252;68mL[38;2;128;255;65mL[38;2;127;255;67mL[38;2;122;255;67mL[38;2;116;255;64mC[38;2;112;251;67mC[38;2;109;238;73mJ[38;2;111;219;79mU[38;2;110;190;91mY[38;2;111;157;103mz[38;2;119;125;126mz[38;2;127;114;140mX[38;2;126;121;137mY[38;2;153;145;152mL[38;2;175;162;171mZ[38;2;134;128;139mU[38;2;124;115;136mX[38;2;101;106;107mn[38;2;78;155;75mn[38;2;71;217;65mc[38;2;72;249;65mY[38;2;71;255;66mY[38;2;66;255;65mY[38;2;63;255;64mX[38;2;58;255;63mX[38;2;58;252;65mX[38;2;60;240;67mz[38;2;63;225;75mz[38;2;75;197;87mz[38;2;94;161;104mz[38;2;112;130;122mz[38;2;126;116;135mX[38;2;132;121;138mY[38;2;109;103;115mu[38;2;33;32;35mI[38;2;0;0;0m   [38;2;0;0;0m");
  $display("[38;2;29;27;26m,[38;2;29;27;25m,[38;2;28;26;24m,[38;2;26;25;23m,[38;2;26;24;24m,[38;2;21;19;19m\"[38;2;29;26;26m,[38;2;56;53;51m~[38;2;103;96;91mx[38;2;150;138;132mJ[38;2;221;204;197ma[38;2;225;206;199ma[38;2;226;207;200mo[38;2;224;207;199ma[38;2;223;207;199ma[38;2;224;207;199maaaa[38;2;227;210;202mo[38;2;218;201;193mh[38;2;168;151;143mQ[38;2;158;139;132mC[38;2;164;145;138mLL[38;2;165;146;139mL[38;2;166;147;140mQ[38;2;156;137;130mJ[38;2;149;130;123mU[38;2;152;133;126mU[38;2;156;136;129mJ[38;2;172;152;145m0[38;2;197;177;170mq[38;2;205;186;179md[38;2;203;184;177md[38;2;193;174;167mw[38;2;181;162;155mZ[38;2;172;153;146m0[38;2;167;148;141mQ[38;2;163;144;137mL[38;2;169;150;143mQ[38;2;220;201;194mh[38;2;226;207;200mo[38;2;225;206;199maa[38;2;222;209;199ma[38;2;232;216;212m#[38;2;167;131;144mL[38;2;77;15;47mi[38;2;83;10;52mi[38;2;84;7;52mi[38;2;82;8;48mi[38;2;80;8;48m!![38;2;81;9;49mi[38;2;82;9;49mi[38;2;94;11;57m~[38;2;111;18;68m-[38;2;113;20;73m-[38;2;103;21;66m_[38;2;126;67;92mr[38;2;171;140;143mQ[38;2;155;136;129mJ[38;2;192;173;167mw[38;2;205;186;179md[38;2;167;148;142mQ[38;2;160;141;135mC[38;2;163;144;137mLLLLLLL[38;2;150;131;124mU[38;2;147;128;121mY[38;2;159;140;133mC[38;2;173;154;147m0[38;2;183;164;155mZ[38;2;162;143;134mC[38;2;158;133;134mJ[38;2;87;36;58m_[38;2;80;9;46m![38;2;82;9;47mi[38;2;79;10;49mi[38;2;81;9;50mi[38;2;81;8;51mi[38;2;82;7;51mi[38;2;83;14;54mi[38;2;124;105;125mc[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;229;79mq[38;2;251;254;72mb[38;2;245;251;71md[38;2;242;252;71md[38;2;241;253;69mp[38;2;243;255;70md[38;2;240;255;71md[38;2;237;255;71mp[38;2;234;255;70mp[38;2;231;255;71mp[38;2;229;255;70mp[38;2;228;255;66mp[38;2;224;255;69mq[38;2;219;255;67mq[38;2;208;249;67mw[38;2;176;209;71mQ[38;2;121;132;84mv[38;2;113;106;121mv[38;2;129;120;142mY[38;2;117;111;125mc[38;2;155;185;85mJ[38;2;195;255;69mm[38;2;188;252;69mZ[38;2;188;254;66mZ[38;2;175;235;72mO[38;2;105;114;95mn[38;2;121;111;133mz[38;2;127;116;145mY[38;2;111;103;125mv[38;2;116;147;84mc[38;2;169;251;71mO[38;2;164;253;68mO[38;2;162;253;66mO[38;2;161;250;72mO[38;2;118;151;93mz[38;2;123;112;138mX[38;2;129;123;137mY[38;2;105;100;109mn[38;2;91;86;94mj[38;2;112;107;117mv[38;2;127;121;136mY[38;2;127;119;140mY[38;2;116;108;129mc[38;2;104;108;107mu[38;2;97;130;84mn[38;2;102;165;75mv[38;2;108;197;71mX[38;2;110;225;65mU[38;2;114;244;66mJ[38;2;116;254;66mC[38;2;113;255;65mC[38;2;108;255;64mC[38;2;106;255;63mJ[38;2;104;254;66mJ[38;2;100;232;72mU[38;2;106;176;94mX[38;2;117;121;124mz[38;2;126;117;135mX[38;2;139;132;145mJ[38;2;146;135;140mJ[38;2;131;122;135mY[38;2;129;120;140mY[38;2;119;110;130mz[38;2;102;108;109mu[38;2;87;125;92mn[38;2;74;159;74mn[38;2;66;194;67mu[38;2;65;219;65mc[38;2;58;243;62mz[38;2;55;255;61mz[38;2;54;255;63mX[38;2;51;255;64mz[38;2;48;255;65mz[38;2;45;255;62mz[38;2;52;237;71mz[38;2;69;190;86mc[38;2;108;127;117mc[38;2;130;121;140mY[38;2;125;118;132mX[38;2;53;48;54m~[38;2;0;0;0m [38;2;0;0;1m [38;2;0;0;1m");
  $display("[38;2;0;0;0m     [38;2;79;73;69m?[38;2;177;162;157mZ[38;2;208;193;186mb[38;2;224;209;201mo[38;2;230;213;206m*[38;2;223;205;198ma[38;2;204;185;178md[38;2;212;193;186mk[38;2;225;208;200mo[38;2;224;207;199maaaaaa[38;2;226;209;201mo[38;2;222;205;197ma[38;2;173;154;147m0[38;2;145;126;120mY[38;2;153;134;127mJ[38;2;155;136;129mJ[38;2;154;135;128mJ[38;2;159;140;133mC[38;2;164;145;138mL[38;2;161;142;135mC[38;2;157;138;131mC[38;2;154;135;128mJ[38;2;154;134;127mJ[38;2;152;133;126mU[38;2;151;132;125mU[38;2;152;133;126mUU[38;2;149;130;123mU[38;2;146;127;120mY[38;2;152;133;126mU[38;2;157;138;131mC[38;2;216;197;190mk[38;2;226;207;200mo[38;2;225;206;199maa[38;2;223;208;199ma[38;2;224;210;202mo[38;2;214;195;195mk[38;2;94;45;66m-[38;2;77;9;48m![38;2;83;8;54mi[38;2;81;8;51mi[38;2;80;8;48m!!!![38;2;83;7;50mi[38;2;97;12;60m+[38;2;112;20;72m-[38;2;113;20;72m-[38;2;105;19;65m_[38;2;132;73;100mn[38;2;159;134;137mC[38;2;166;150;143mQ[38;2;226;207;201mo[38;2;218;198;193mh[38;2;182;163;156mZ[38;2;160;141;134mC[38;2;161;142;135mC[38;2;162;143;136mL[38;2;163;144;137mLLL[38;2;159;140;132mC[38;2;152;133;126mU[38;2;186;167;160mm[38;2;183;164;157mZ[38;2;223;204;197ma[38;2;228;207;199mo[38;2;191;174;165mw[38;2;163;143;142mL[38;2;101;56;75m1[38;2;78;8;45m![38;2;82;10;49mi[38;2;78;9;48m![38;2;79;7;49m![38;2;80;7;50m![38;2;81;6;49m![38;2;86;17;57m~[38;2;125;107;127mz[38;2;127;122;140mY[38;2;114;113;103mv[38;2;230;229;79mq[38;2;251;254;72mb[38;2;245;251;71md[38;2;243;253;71md[38;2;234;245;71mp[38;2;205;215;66mO[38;2;202;216;69mO[38;2;200;216;69mO[38;2;197;216;67mO[38;2;195;215;67m0[38;2;189;213;72m0[38;2;180;203;73mQ[38;2;165;183;74mJ[38;2;142;155;78mX[38;2;119;124;90mv[38;2;107;106;113mu[38;2;119;113;135mz[38;2;130;121;141mY[38;2;122;115;130mz[38;2;130;148;95mX[38;2;195;249;72mm[38;2;190;254;66mm[38;2;189;252;69mm[38;2;189;255;67mm[38;2;159;210;73mL[38;2;130;153;88mz[38;2;141;166;105mU[38;2;138;166;101mU[38;2;139;164;104mU[38;2;121;158;82mz[38;2;159;236;70mQ[38;2;165;254;69mO[38;2;162;252;68mO[38;2;162;255;66mO[38;2;148;228;74mL[38;2;112;122;110mv[38;2;129;118;137mY[38;2;122;119;133mX[38;2;123;116;132mz[38;2;128;118;137mX[38;2;124;116;135mX[38;2;126;116;137mX[38;2;128;117;135mX[38;2;125;116;140mX[38;2;127;113;138mX[38;2;120;109;130mz[38;2;112;105;121mv[38;2;104;108;108mu[38;2;99;119;95mn[38;2;93;138;82mn[38;2;93;171;70mv[38;2;100;217;66mX[38;2;107;253;68mC[38;2;103;253;65mJ[38;2;101;254;67mJ[38;2;99;255;68mJ[38;2;95;210;74mX[38;2;110;121;117mc[38;2;130;117;138mY[38;2;127;120;137mY[38;2;128;117;137mX[38;2;128;116;138mX[38;2;129;116;139mY[38;2;129;116;140mY[38;2;130;113;141mY[38;2;123;110;133mz[38;2;113;106;122mv[38;2;102;108;111mu[38;2;91;116;99mn[38;2;78;133;83mx[38;2;63;164;72mx[38;2;55;207;68mv[38;2;49;250;62mz[38;2;49;253;67mz[38;2;44;255;62mz[38;2;37;255;59mc[38;2;52;225;74mc[38;2;97;130;109mv[38;2;131;120;142mY[38;2;125;119;132mX[38;2;27;25;28m,[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;0;0;0m    [38;2;16;13;12m'[38;2;197;183;176mp[38;2;236;217;209m#[38;2;227;209;202mo[38;2;225;207;199ma[38;2;224;207;199maa[38;2;224;205;198ma[38;2;207;188;181mb[38;2;201;182;175mp[38;2;224;205;198ma[38;2;225;208;200mo[38;2;224;207;199maaaaa[38;2;225;208;200mo[38;2;226;207;201mo[38;2;180;161;155mZ[38;2;154;135;129mJ[38;2;159;140;134mC[38;2;158;139;132mC[38;2;160;141;134mC[38;2;162;143;136mL[38;2;163;144;137mLLLL[38;2;164;145;138mL[38;2;161;142;135mC[38;2;155;136;129mJ[38;2;151;132;125mU[38;2;149;130;123mUU[38;2;161;141;134mC[38;2;164;145;138mL[38;2;212;193;186mk[38;2;227;208;201mo[38;2;226;207;200mo[38;2;225;206;198ma[38;2;224;207;197ma[38;2;224;207;199ma[38;2;228;212;204mo[38;2;133;98;107mv[38;2;70;13;43m![38;2;81;9;51mi[38;2;82;9;48mi[38;2;82;7;48m![38;2;81;8;48m![38;2;80;8;48m![38;2;79;8;48m![38;2;81;8;49mi[38;2;85;6;51mi[38;2;96;12;60m+[38;2;111;21;72m-[38;2;115;19;73m?[38;2;103;20;66m_[38;2;128;76;101mn[38;2;160;137;138mC[38;2;185;166;163mm[38;2;226;208;202mo[38;2;225;207;200ma[38;2;200;181;175mp[38;2;169;150;143mQ[38;2;159;141;131mC[38;2;161;143;133mCC[38;2;164;146;136mL[38;2;184;166;156mZ[38;2;212;193;186mk[38;2;217;198;191mh[38;2;196;177;170mq[38;2;228;208;201mo[38;2;226;207;198ma[38;2;224;209;199ma[38;2;197;177;174mq[38;2;120;86;99mn[38;2;73;11;45m![38;2;80;11;51mi[38;2;79;10;49mi[38;2;80;8;47m![38;2;80;8;49m![38;2;84;5;50mi[38;2;97;22;66m_[38;2;127;108;128mz[38;2;125;123;140mY[38;2;117;111;103mv[38;2;229;230;78mq[38;2;251;255;71mb[38;2;245;252;71md[38;2;246;255;72md[38;2;209;220;74mZ[38;2;102;96;94mx[38;2;109;106;116mv[38;2;111;106;115mv[38;2;112;107;113mv[38;2;112;107;115mv[38;2;112;106;116mv[38;2;112;106;120mv[38;2;115;107;128mc[38;2;120;111;134mz[38;2;124;116;136mX[38;2;126;119;135mX[38;2;129;122;141mY[38;2;125;120;138mX[38;2;117;120;111mc[38;2;183;226;78mO[38;2;198;255;69mw[38;2;192;253;66mm[38;2;188;253;71mm[38;2;189;255;68mmm[38;2;189;255;67mm[38;2;185;255;67mZ[38;2;180;255;68mZ[38;2;177;255;68mZ[38;2;174;255;68mZ[38;2;168;255;69mO[38;2;164;255;68mO[38;2;161;253;67mO[38;2;159;252;69mO[38;2;158;255;71mO[38;2;135;193;79mU[38;2;115;111;126mc[38;2;129;121;142mY[38;2;125;115;133mX[38;2;121;152;106mX[38;2;130;204;90mJ[38;2;128;200;90mJ[38;2;128;200;88mJ[38;2;127;201;91mJ[38;2;119;144;105mz[38;2;126;114;139mX[38;2;130;122;139mY[38;2;131;122;140mY[38;2;128;119;139mY[38;2;128;113;137mX[38;2;114;109;128mc[38;2;97;98;104mx[38;2;93;185;71mc[38;2;105;255;68mC[38;2;99;253;67mJ[38;2;97;254;65mJ[38;2;98;255;67mJ[38;2;92;153;88mv[38;2;127;107;137mz[38;2;106;139;111mc[38;2;97;201;93mY[38;2;94;200;89mXX[38;2;91;202;87mX[38;2;101;159;101mz[38;2;123;114;136mX[38;2;130;123;138mY[38;2;129;121;139mY[38;2;129;118;138mY[38;2;128;115;138mX[38;2;122;108;132mz[38;2;104;97;111mn[38;2;62;159;73mx[38;2;50;253;66mz[38;2;44;254;66mz[38;2;42;254;63mz[38;2;36;255;65mc[38;2;63;178;78mu[38;2;119;111;133mz[38;2;134;127;143mU[38;2;68;65;73m-[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;0;0;0m    [38;2;15;11;10m'[38;2;190;175;169mw[38;2;229;210;203mo[38;2;224;207;199maaaa[38;2;225;206;199ma[38;2;227;208;201mo[38;2;216;197;190mk[38;2;198;179;172mp[38;2;218;201;193mh[38;2;226;209;201mo[38;2;224;207;199maaaaa[38;2;226;207;201mo[38;2;229;210;204mo[38;2;189;170;164mw[38;2;158;139;133mC[38;2;163;144;137mL[38;2;162;143;136mLLLL[38;2;163;144;137mL[38;2;161;142;135mC[38;2;152;132;125mU[38;2;147;127;120mY[38;2;150;131;124mU[38;2;158;139;132mC[38;2;166;148;140mQ[38;2;173;155;147m0[38;2;172;153;146m0[38;2;172;154;146m0[38;2;199;180;173mp[38;2;216;197;190mk[38;2;223;204;197ma[38;2;226;208;200mo[38;2;224;207;197ma[38;2;224;207;199ma[38;2;228;212;204mo[38;2;179;161;156mZ[38;2;124;93;97mn[38;2;83;32;54m+[38;2;75;8;43m![38;2;83;8;49mi[38;2;82;8;49mi[38;2;80;8;48m![38;2;79;8;48m![38;2;81;8;48m![38;2;82;7;50mi[38;2;84;7;52mi[38;2;94;15;61m+[38;2;112;20;72m-[38;2;115;18;72m-[38;2;104;23;66m-[38;2;129;84;102mn[38;2;178;157;158mO[38;2;196;183;175mp[38;2;223;205;198ma[38;2;228;209;203mo[38;2;219;200;193mh[38;2;193;175;165mw[38;2;177;159;149mO[38;2;188;170;161mm[38;2;211;193;183mb[38;2;226;208;198ma[38;2;227;208;200mo[38;2;222;203;196ma[38;2;190;172;165mw[38;2;224;206;199ma[38;2;224;208;199ma[38;2;222;209;197ma[38;2;227;210;205mo[38;2;168;142;149mQ[38;2;75;22;49mi[38;2;82;10;51mi[38;2;79;10;53mi[38;2;78;9;49m![38;2;80;7;48m![38;2;92;8;55m~[38;2;107;24;71m-[38;2;127;107;128mz[38;2;124;123;140mY[38;2;117;111;103mv[38;2;229;230;78mq[38;2;251;255;71mb[38;2;245;251;70md[38;2;245;255;71md[38;2;209;219;76mZ[38;2;115;108;114mv[38;2;127;122;141mY[38;2;127;120;137mY[38;2;118;110;126mc[38;2;116;109;124mc[38;2;123;116;130mz[38;2;125;119;131mX[38;2;120;114;123mz[38;2;104;98;107mn[38;2;98;93;101mx[38;2;120;113;126mz[38;2;131;121;140mY[38;2;116;112;121mc[38;2;159;190;88mC[38;2;202;255;66mw[38;2;195;252;66mm[38;2;192;253;69mm[38;2;188;250;71mZ[38;2;158;208;66mC[38;2;154;204;68mC[38;2;153;205;69mC[38;2;151;204;70mJ[38;2;149;204;69mJ[38;2;146;205;68mJ[38;2;144;205;67mJ[38;2;139;202;70mU[38;2;147;220;67mC[38;2;164;254;70mO[38;2;157;253;68m0[38;2;157;253;67m0[38;2;155;251;68m0[38;2;120;154;93mz[38;2;123;112;136mz[38;2;124;114;136mX[38;2;104;137;86mu[38;2;143;254;67mQ[38;2;137;255;65mQ[38;2;137;255;68mQ[38;2;131;255;63mL[38;2;122;211;74mU[38;2;112;125;115mc[38;2;124;115;134mX[38;2;129;114;140mX[38;2;128;116;137mX[38;2;130;114;141mY[38;2;127;116;139mX[38;2;117;111;123mc[38;2;97;184;77mz[38;2;104;255;68mC[38;2;100;253;68mJ[38;2;96;254;64mJ[38;2;96;255;67mJ[38;2;90;149;87mu[38;2;125;108;132mz[38;2;94;120;97mn[38;2;84;238;70mY[38;2;79;255;64mY[38;2;77;255;65mY[38;2;72;255;62mY[38;2;73;231;71mX[38;2;100;135;101mv[38;2;124;115;137mX[38;2;127;115;137mX[38;2;128;115;139mX[38;2;130;115;140mY[38;2;129;116;138mX[38;2;122;113;129mz[38;2;73;160;87mu[38;2;50;253;65mz[38;2;44;254;66mz[38;2;42;253;63mz[38;2;35;255;63mc[38;2;62;176;75mn[38;2;114;109;129mc[38;2;134;127;144mU[38;2;71;68;75m?[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;0;0;0m    [38;2;3;1;1m [38;2;157;144;141mL[38;2;233;216;208m*[38;2;225;208;199ma[38;2;225;208;200mooooo[38;2;227;210;202mo[38;2;220;203;195ma[38;2;199;182;174mp[38;2;211;194;186mk[38;2;225;208;200mo[38;2;224;207;199maaa[38;2;225;208;200mo[38;2;227;209;202mo[38;2;216;197;191mk[38;2;204;185;179md[38;2;165;146;140mL[38;2;154;135;128mJ[38;2;163;144;137mL[38;2;162;143;136mLL[38;2;163;144;137mL[38;2;154;135;128mJ[38;2;144;125;118mY[38;2;157;137;130mJ[38;2;179;160;153mO[38;2;199;180;173mp[38;2;212;193;186mk[38;2;216;199;191mh[38;2;222;205;197ma[38;2;225;208;200moo[38;2;223;206;198ma[38;2;222;205;197ma[38;2;224;207;199maaaa[38;2;227;210;202mo[38;2;198;179;170mq[38;2;155;136;123mJ[38;2;154;128;126mU[38;2;98;57;77m1[38;2;74;13;47m![38;2;80;8;50mi[38;2;83;7;50mi[38;2;81;8;48m![38;2;80;7;50m![38;2;81;8;51mii[38;2;83;9;51mi[38;2;93;11;57m~[38;2;107;17;67m_[38;2;111;19;72m-[38;2;100;25;69m-[38;2;140;101;116mz[38;2;203;185;179md[38;2;221;201;195mh[38;2;225;206;200ma[38;2;226;207;200mo[38;2;227;208;201mo[38;2;225;206;199ma[38;2;227;208;201moo[38;2;225;206;199ma[38;2;224;207;199ma[38;2;226;209;201mo[38;2;200;183;175mp[38;2;207;191;184mb[38;2;227;208;202mo[38;2;224;207;196ma[38;2;230;213;207m*[38;2;194;154;149mZ[38;2;94;34;46m+[38;2;83;9;48mi[38;2;81;9;51mi[38;2;79;9;49m![38;2;83;8;50mi[38;2;100;14;61m+[38;2;109;25;72m-[38;2;127;107;128mz[38;2;124;123;140mY[38;2;117;111;103mv[38;2;229;230;78mq[38;2;251;255;71mb[38;2;245;251;70md[38;2;245;255;71md[38;2;209;220;76mZ[38;2;114;108;111mv[38;2;126;122;140mY[38;2;122;115;131mz[38;2;104;95;105mn[38;2;110;103;113mu[38;2;117;111;121mc[38;2;116;112;120mc[38;2;120;113;119mc[38;2;116;109;115mv[38;2;114;106;119mv[38;2;129;121;137mY[38;2;120;114;136mz[38;2;135;150;95mX[38;2;202;250;72mw[38;2;197;254;68mm[38;2;196;252;66mm[38;2;194;255;69mm[38;2;153;193;73mJ[38;2;99;95;102mx[38;2;112;106;119mv[38;2;115;109;123mc[38;2;118;112;125mcc[38;2;118;111;126mc[38;2;116;110;124mc[38;2;110;103;120mv[38;2;95;109;89mx[38;2;151;229;71mL[38;2;160;255;67mO[38;2;158;252;68m0[38;2;154;255;68m0[38;2;149;231;69mL[38;2;112;124;111mc[38;2;130;117;141mY[38;2;113;105;122mv[38;2;103;155;77mv[38;2;135;242;68mL[38;2;136;255;68mQ[38;2;131;255;66mL[38;2;130;255;65mL[38;2;125;238;69mC[38;2;118;206;82mU[38;2;117;185;97mU[38;2;114;179;96mY[38;2;113;178;98mY[38;2;114;189;92mY[38;2;109;219;75mU[38;2;107;251;69mC[38;2;106;252;68mC[38;2;100;255;64mJ[38;2;98;255;66mJ[38;2;91;206;72mz[38;2;101;110;105mn[38;2;130;118;140mY[38;2;115;111;126mc[38;2;84;134;84mx[38;2;78;231;69mX[38;2;78;255;67mU[38;2;75;255;65mY[38;2;69;255;64mY[38;2;73;244;68mY[38;2;80;210;82mX[38;2;86;188;92mz[38;2;89;178;95mz[38;2;87;178;95mz[38;2;84;187;90mz[38;2;70;211;80mz[38;2;49;249;68mz[38;2;48;254;66mz[38;2;44;255;68mz[38;2;42;255;62mz[38;2;40;226;66mv[38;2;84;119;94mx[38;2;128;117;137mX[38;2;129;122;138mY[38;2;34;33;37mI[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;0;0;0m     [38;2;80;74;71m1[38;2;215;200;195mh[38;2;229;211;204mo[38;2;227;210;203mo[38;2;226;209;201mo[38;2;225;208;200moooo[38;2;226;209;201moo[38;2;207;190;182mb[38;2;206;189;181mb[38;2;225;208;200moo[38;2;227;210;202mo[38;2;223;206;198ma[38;2;196;178;171mq[38;2;168;149;143mQ[38;2;160;141;135mC[38;2;157;138;132mC[38;2;146;127;120mY[38;2;163;144;137mLL[38;2;161;142;135mC[38;2;146;127;120mY[38;2;152;133;126mU[38;2;188;169;162mm[38;2;215;197;190mk[38;2;225;208;200mo[38;2;228;211;203mo[38;2;226;209;201mo[38;2;225;208;200moo[38;2;224;207;199maaaaaaaa[38;2;226;209;202mo[38;2;212;188;178mb[38;2;155;101;79mv[38;2;177;106;84mz[38;2;173;115;104mY[38;2;126;75;76mr[38;2;81;18;42mi[38;2;77;7;47m![38;2;80;9;52mi[38;2;80;7;50m![38;2;80;7;49m![38;2;80;7;50m![38;2;82;9;51mi[38;2;82;8;51mi[38;2;89;10;56m~[38;2;106;18;69m-[38;2;111;19;71m-[38;2;102;31;73m-[38;2;167;128;144mC[38;2;225;207;200ma[38;2;226;207;199ma[38;2;225;206;199maaaaaa[38;2;224;207;199maa[38;2;223;206;198ma[38;2;195;177;170mq[38;2;220;201;194mh[38;2;229;213;206m*[38;2;209;168;159mw[38;2;182;97;70mc[38;2;144;54;45mt[38;2;84;8;41m![38;2;80;9;49mi[38;2;82;9;47mi[38;2;88;9;52mi[38;2;106;17;65m_[38;2;112;24;74m?[38;2;127;108;129mz[38;2;124;123;139mY[38;2;117;111;101mu[38;2;232;235;78mq[38;2;255;255;71mb[38;2;250;255;70md[38;2;251;255;71mb[38;2;213;224;75mm[38;2;113;108;110mv[38;2;126;122;139mY[38;2;125;118;135mX[38;2;115;109;119mv[38;2;116;112;121mc[38;2;114;113;121mc[38;2;115;113;121mc[38;2;119;111;122mc[38;2;121;114;124mz[38;2;130;121;137mY[38;2;127;117;140mY[38;2;122;126;106mc[38;2;194;236;76mZ[38;2;208;255;65mw[38;2;201;255;67mw[38;2;200;255;65mm[38;2;184;239;70mO[38;2;108;116;92mn[38;2;123;116;137mX[38;2;130;124;138mY[38;2;86;80;89mf[38;2;62;58;66m_[38;2;65;61;68m-[38;2;64;60;68m-[38;2;90;84;98mj[38;2;132;126;141mU[38;2;117;107;130mc[38;2;111;148;77mv[38;2;163;255;71mO[38;2;158;255;67mO[38;2;155;255;66m0[38;2;153;255;65m0[38;2;134;203;81mJ[38;2;116;115;121mc[38;2;131;119;137mY[38;2;114;107;128mc[38;2;99;121;87mn[38;2;113;176;76mz[38;2;121;226;65mU[38;2;126;250;63mC[38;2;128;255;67mL[38;2;125;255;64mL[38;2;121;255;62mC[38;2;120;255;65mC[38;2;115;255;64mC[38;2;113;255;64mC[38;2;110;255;65mC[38;2;105;255;65mJ[38;2;102;249;67mJ[38;2;95;222;63mX[38;2;89;162;75mu[38;2;97;109;104mn[38;2;126;116;137mX[38;2;127;122;136mY[38;2;127;122;137mY[38;2;121;109;132mz[38;2;94;112;100mn[38;2;74;168;71mn[38;2;72;220;65mz[38;2;73;246;64mX[38;2;69;255;64mY[38;2;64;255;63mX[38;2;62;255;63mX[38;2;60;255;63mX[38;2;57;255;62mX[38;2;53;255;61mz[38;2;50;255;62mz[38;2;47;255;67mz[38;2;46;252;61mz[38;2;46;231;64mv[38;2;55;177;70mx[38;2;88;114;95mx[38;2;127;114;136mX[38;2;131;126;140mY[38;2;67;63;70m-[38;2;1;0;1m [38;2;0;0;0m [38;2;0;0;1m");
  $display("[38;2;0;0;0m   [38;2;43;42;41m![38;2;131;130;127mY[38;2;158;150;148mQ[38;2;154;137;136mC[38;2;182;163;161mZ[38;2;209;191;187mb[38;2;224;206;201ma[38;2;228;211;204mo[38;2;226;207;200moo[38;2;228;209;202mo[38;2;229;210;203mo[38;2;224;206;199ma[38;2;217;198;191mh[38;2;194;175;168mq[38;2;186;168;160mm[38;2;220;203;195ma[38;2;209;192;184mb[38;2;172;155;147m0[38;2;153;134;127mJ[38;2;150;131;124mU[38;2;143;124;117mY[38;2;147;128;121mY[38;2;144;125;118mY[38;2;164;145;138mL[38;2;159;140;133mC[38;2;143;124;117mY[38;2;167;148;141mQ[38;2;212;193;186mk[38;2;228;209;202mo[38;2;226;209;201mo[38;2;224;207;199maaaaaaaaaaaaa[38;2;225;209;201mo[38;2;216;196;185mk[38;2;176;104;70mc[38;2;204;90;41mv[38;2;199;90;46mv[38;2;195;93;54mv[38;2;169;72;52mx[38;2;108;25;39m+[38;2;77;6;43m![38;2;80;9;50mi[38;2;83;8;47mi[38;2;81;7;47m![38;2;78;8;48m![38;2;79;8;49m![38;2;82;7;50mi[38;2;87;9;55mi[38;2;102;17;66m_[38;2;107;18;69m-[38;2;111;50;79mt[38;2;194;168;169mw[38;2;227;210;203mo[38;2;224;207;196ma[38;2;224;207;198ma[38;2;224;207;200ma[38;2;224;207;199maaaa[38;2;222;208;199ma[38;2;225;208;200mo[38;2;224;205;198ma[38;2;225;205;198ma[38;2;204;159;146mZ[38;2;184;96;69mc[38;2;206;93;48mc[38;2;182;80;51mn[38;2;94;14;33mi[38;2;80;8;49m![38;2;82;7;49mi[38;2;89;8;53mi[38;2;107;17;67m_[38;2;111;21;72m-[38;2;127;100;122mc[38;2;125;123;141mY[38;2;118;111;113mv[38;2;147;147;89mX[38;2;151;154;80mY[38;2;150;152;80mX[38;2;151;153;79mX[38;2;142;144;88mX[38;2;118;112;126mc[38;2;128;122;138mY[38;2;125;118;136mX[38;2;116;113;119mc[38;2;116;113;122mc[38;2;115;112;121mcc[38;2;117;111;123mc[38;2;122;115;129mz[38;2;128;121;137mY[38;2;123;116;138mX[38;2;123;129;101mc[38;2;138;156;82mX[38;2;134;152;83mz[38;2;132;152;79mz[38;2;130;156;78mz[38;2;121;136;91mc[38;2;117;111;126mc[38;2;126;120;138mY[38;2;148;141;145mC[38;2;133;128;114mX[38;2;14;12;8m'[38;2;0;0;0m  [38;2;10;9;12m'[38;2;108;104;112mu[38;2;136;125;147mU[38;2;111;112;117mv[38;2;116;148;87mc[38;2;114;155;79mc[38;2;113;153;80mc[38;2;110;152;79mv[38;2;115;152;84mc[38;2;110;121;110mv[38;2;124;117;138mX[38;2;130;120;135mY[38;2;124;115;139mX[38;2;111;103;122mv[38;2;103;106;105mn[38;2;98;125;88mn[38;2;97;149;81mu[38;2;102;165;77mv[38;2;102;173;71mc[38;2;99;176;72mc[38;2;95;177;72mv[38;2;97;174;69mv[38;2;95;165;76mv[38;2;92;149;82mu[38;2;95;125;89mn[38;2;103;107;108mu[38;2;117;108;128mc[38;2;127;120;138mY[38;2;128;118;127mX[38;2;131;117;117mz[38;2;138;125;125mY[38;2;131;122;134mY[38;2;129;118;139mY[38;2;118;107;130mc[38;2;101;107;110mu[38;2;89;120;94mn[38;2;77;143;81mx[38;2;71;164;75mn[38;2;68;172;73mn[38;2;66;175;72mn[38;2;65;176;72mn[38;2;64;175;71mn[38;2;62;168;74mn[38;2;67;154;78mx[38;2;80;131;88mx[38;2;98;113;107mu[38;2;121;111;131mz[38;2;132;122;142mY[38;2;111;105;116mv[38;2;48;45;52mi[38;2;0;0;0m   [38;2;0;0;0m");
  $display("[38;2;69;67;65m-[38;2;118;115;113mc[38;2;179;176;174mw[38;2;230;229;226mM[38;2;247;248;244mB[38;2;215;209;206ma[38;2;150;138;135mJ[38;2;149;133;131mU[38;2;147;129;126mU[38;2;156;138;133mC[38;2;199;182;175mp[38;2;226;208;201mo[38;2;227;208;201mo[38;2;216;197;190mk[38;2;194;174;167mw[38;2;174;155;147m0[38;2;165;146;139mL[38;2;164;145;138mL[38;2;160;142;134mC[38;2;154;137;129mJ[38;2;163;145;137mL[38;2;159;142;134mC[38;2;157;138;131mC[38;2;156;137;130mJ[38;2;149;130;123mU[38;2;160;141;134mC[38;2;143;124;117mY[38;2;161;142;135mC[38;2;142;123;116mX[38;2;168;149;142mQ[38;2;219;200;193mh[38;2;229;210;203mo[38;2;226;207;200mo[38;2;225;208;200moooooooooooooo[38;2;226;210;202mo[38;2;215;196;186mk[38;2;166;107;86mz[38;2;193;96;62mc[38;2;194;91;51mv[38;2;201;91;46mv[38;2;210;94;48mc[38;2;192;87;55mv[38;2;132;44;38m?[38;2;86;12;38m![38;2;80;9;51mi[38;2;81;9;48mi[38;2;81;8;46m![38;2;81;7;49m![38;2;81;7;50mi[38;2;82;8;52mi[38;2;86;9;53mi[38;2;104;13;66m_[38;2;103;20;67m_[38;2;137;83;105mu[38;2;217;189;185mk[38;2;232;210;198mo[38;2;228;211;202mo[38;2;227;211;203mo[38;2;226;209;201mo[38;2;225;208;200moo[38;2;225;208;199ma[38;2;223;209;200ma[38;2;227;211;203mo[38;2;225;198;189mh[38;2;195;137;119mL[38;2;189;91;54mv[38;2;206;91;46mv[38;2;201;93;49mv[38;2;184;104;78mz[38;2;128;76;88mx[38;2;75;10;47m![38;2;82;8;50mi[38;2;87;9;53mi[38;2;105;18;67m_[38;2;112;18;71m-[38;2;113;39;83mt[38;2;137;116;136mY[38;2;141;135;148mJ[38;2;124;118;140mX[38;2;121;116;138mX[38;2;122;117;138mXX[38;2;125;118;141mY[38;2;127;121;136mY[38;2;125;119;129mX[38;2;119;114;124mz[38;2;115;113;121mc[38;2;115;113;122mc[38;2;116;112;121mcc[38;2;118;112;120mc[38;2;118;112;123mc[38;2;123;117;129mz[38;2;125;121;134mX[38;2;124;117;136mX[38;2;122;111;136mz[38;2;120;112;135mz[38;2;120;112;133mz[38;2;121;112;134mz[38;2;123;115;135mX[38;2;125;118;133mX[38;2;145;143;146mC[38;2;168;171;155mO[38;2;180;180;166mw[38;2;108;106;94mn[38;2;3;3;2m [38;2;0;0;1m [38;2;0;0;0m [38;2;23;20;24m\"[38;2;87;85;93mj[38;2;115;111;126mc[38;2;121;110;132mz[38;2;119;109;132mz[38;2;119;110;133mz[38;2;125;115;138mX[38;2;126;116;138mX[38;2;134;126;142mU[38;2;151;140;149mC[38;2;189;177;178mq[38;2;195;182;182mp[38;2;167;156;162mO[38;2;147;138;151mC[38;2;131;120;140mY[38;2;126;113;137mX[38;2;122;110;132mz[38;2;120;108;130mz[38;2;121;108;131mz[38;2;121;108;132mz[38;2;121;109;131mz[38;2;121;111;132mz[38;2;124;113;136mX[38;2;127;116;138mX[38;2;135;125;139mU[38;2;135;123;131mY[38;2;155;139;141mC[38;2;159;140;135mC[38;2;146;126;116mY[38;2;152;135;125mU[38;2;159;141;136mC[38;2;153;137;135mJ[38;2;143;132;136mU[38;2;137;126;140mU[38;2;134;121;141mY[38;2;130;117;136mX[38;2;124;112;130mz[38;2;120;109;128mz[38;2;119;109;129mz[38;2;120;108;129mz[38;2;123;109;131mz[38;2;125;110;134mz[38;2;125;112;135mX[38;2;123;111;132mz[38;2;110;102;120mv[38;2;83;80;92mf[38;2;44;43;50m![38;2;8;8;8m.[38;2;0;0;0m    [38;2;0;0;0m");
  $display("[38;2;226;226;226mM[38;2;233;233;231mW[38;2;231;231;227mW[38;2;226;227;222mM[38;2;224;225;221m#[38;2;229;227;223mM[38;2;179;173;170mw[38;2;143;132;130mU[38;2;152;138;133mJ[38;2;151;136;130mJ[38;2;147;130;123mU[38;2;152;134;128mJ[38;2;172;153;147m0[38;2;162;142;134mC[38;2;156;134;126mJ[38;2;157;137;129mJ[38;2;156;139;129mJ[38;2;154;138;129mJ[38;2;155;139;130mJ[38;2;142;124;117mX[38;2;140;122;114mX[38;2;158;140;132mC[38;2;155;138;130mJ[38;2;154;137;130mJ[38;2;155;139;131mJ[38;2;155;138;130mJ[38;2;132;114;107mc[38;2;149;131;124mU[38;2;148;130;122mU[38;2;194;177;169mq[38;2;217;200;192mh[38;2;215;198;190mk[38;2;214;197;190mkkkkkkkkkkkkkkk[38;2;215;199;191mk[38;2;201;186;181md[38;2;190;175;168mw[38;2;210;190;180mb[38;2;190;161;148mZ[38;2;183;130;114mC[38;2;177;101;78mc[38;2;176;90;58mu[38;2;188;89;60mv[38;2;139;52;46mt[38;2;80;11;39m![38;2;77;10;45m![38;2;78;9;45m![38;2;76;7;46m![38;2;77;8;46m![38;2;77;8;47m![38;2;75;8;46m![38;2;82;9;50mi[38;2;97;18;64m+[38;2;101;23;61m_[38;2;153;89;84mu[38;2;186;131;106mJ[38;2;195;152;136mO[38;2;206;174;162mq[38;2;215;193;184mk[38;2;214;198;191mk[38;2;213;198;188mk[38;2;215;198;188mk[38;2;217;199;194mh[38;2;201;177;164mq[38;2;172;110;87mz[38;2;183;82;49mn[38;2;196;87;46mu[38;2;192;87;47mu[38;2;174;93;64mv[38;2;209;185;173md[38;2;196;188;193mb[38;2;77;26;54m~[38;2;75;8;46m![38;2;81;8;48m![38;2;98;15;61m+[38;2;107;19;69m-[38;2;97;14;60m+[38;2;160;125;144mC[38;2;221;218;222m#[38;2;202;202;203mhhh[38;2;203;203;204mh[38;2;206;206;208ma[38;2;153;152;155mQ[38;2;106;105;104mn[38;2;109;109;113mv[38;2;109;108;117mv[38;2;109;107;116mv[38;2;111;106;116mv[38;2;112;106;116mv[38;2;113;107;117mvv[38;2;112;106;116mv[38;2;111;106;117mv[38;2;112;108;119mv[38;2;113;109;119mv[38;2;113;110;121mv[38;2;106;103;114mu[38;2;91;87;96mj[38;2;95;92;99mr[38;2;92;90;95mr[38;2;138;139;133mU[38;2;163;167;151mOO[38;2;154;154;141mL[38;2;28;25;22m,[38;2;0;0;0m [38;2;0;0;2m [38;2;0;0;0m  [38;2;13;13;14m'[38;2;25;26;27m,[38;2;26;25;29m,[38;2;37;33;36mI[38;2;166;155;155m0[38;2;198;183;180mp[38;2;202;186;181md[38;2;213;197;191mk[38;2;217;201;194mh[38;2;217;201;192mh[38;2;218;202;195mh[38;2;192;174;171mq[38;2;153;137;134mJ[38;2;145;133;133mU[38;2;143;132;133mU[38;2;144;132;135mU[38;2;126;114;118mz[38;2;101;93;100mx[38;2;101;97;104mx[38;2;98;97;104mx[38;2;95;93;101mx[38;2;104;94;99mx[38;2;146;128;125mU[38;2;138;119;111mz[38;2;159;141;132mC[38;2;158;140;132mC[38;2;148;130;123mU[38;2;151;134;126mU[38;2;156;137;130mJ[38;2;156;137;129mJ[38;2;155;137;129mJ[38;2;160;143;136mC[38;2;191;175;170mw[38;2;195;182;178mp[38;2;186;171;172mw[38;2;181;169;172mw[38;2;181;169;169mm[38;2;185;172;172mw[38;2;139;131;135mU[38;2;44;42;49m![38;2;35;33;38mI[38;2;22;21;24m\"[38;2;6;6;9m.[38;2;0;0;0m       [38;2;0;0;0m");
  $display("");
  $display("\033[1;0m");
  $display ("--------------------------------------------------");
  $display("                  Congratulations!               ");
  $display("              execution cycles = %7d", total_latency);
  $display("              clock period = %4fns", CYCLE);
  $display ("--------------------------------------------------");
  $finish;	
endtask

task fail_task;
  $display("[38;2;0;0;0m                                                                   [38;2;2;1;2m [38;2;2;1;3m [38;2;7;5;6m.[38;2;7;5;5m.[38;2;6;4;5m.[38;2;10;9;7m.[38;2;16;14;13m^[38;2;14;12;11m'[38;2;24;23;15m\"[38;2;23;22;15m\"[38;2;28;26;18m,[38;2;38;35;24mI[38;2;40;39;23mI[38;2;50;51;29m![38;2;53;54;30m![38;2;52;50;26m![38;2;59;57;31mi[38;2;82;80;55m?[38;2;91;91;69mf[38;2;55;55;42mi[38;2;29;29;18m,[38;2;73;74;49m-[38;2;63;63;50m+[38;2;4;4;4m [38;2;0;0;0m                                                                                   [38;2;0;0;0m");
  $display("[38;2;0;0;0m                                           [38;2;0;0;2m  [38;2;0;0;1m [38;2;1;0;1m [38;2;6;5;5m.[38;2;10;9;7m.[38;2;9;8;5m.[38;2;11;11;9m'[38;2;11;9;9m.[38;2;23;21;18m\"[38;2;27;25;16m\"[38;2;29;24;17m,[38;2;37;28;18m,[38;2;43;34;20mI[38;2;34;26;16m,[38;2;40;36;20mI[38;2;71;70;40m_[38;2;65;60;32m~[38;2;51;47;26ml[38;2;69;69;48m_[38;2;78;83;57m?[38;2;80;89;56m1[38;2;114;121;98mv[38;2;86;94;84mj[38;2;37;44;30ml[38;2;82;82;60m1[38;2;64;63;40m+[38;2;85;91;51m1[38;2;117;125;73mn[38;2;118;123;74mn[38;2;110;109;60mr[38;2;135;124;67mu[38;2;151;131;65mc[38;2;145;125;54mu[38;2;168;149;69mY[38;2;193;175;85mQ[38;2;189;176;77mL[38;2;170;162;77mU[38;2;192;186;94m0[38;2;208;197;89mO[38;2;200;186;82m0[38;2;190;182;95mQ[38;2;221;219;154mk[38;2;164;160;114mC[38;2;111;106;65mr[38;2;144;140;88mX[38;2;79;75;57m?[38;2;1;1;1m [38;2;0;0;0m                                                                                   [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;2;2;2m [38;2;14;14;11m'[38;2;11;10;6m.[38;2;23;21;14m\"[38;2;34;30;22m;[38;2;27;22;14m\"[38;2;24;20;14m\"[38;2;36;33;22m;[38;2;51;47;28m![38;2;58;54;28mi[38;2;66;61;31m~[38;2;71;65;34m+[38;2;69;62;30m~[38;2;82;73;35m_[38;2;95;87;41m1[38;2;104;93;46mt[38;2;115;105;54mj[38;2;114;103;45mj[38;2;137;128;62mu[38;2;163;156;89mU[38;2;164;157;93mJ[38;2;143;135;74mc[38;2;133;123;62mu[38;2;114;105;47mj[38;2;126;118;67mn[38;2;154;143;106mU[38;2;175;161;109mL[38;2;186;175;87mL[38;2;138;119;60mn[38;2;133;96;51mr[38;2;207;164;80mL[38;2;184;142;68mY[38;2;137;110;38mr[38;2;198;186;83mQ[38;2;220;207;97mw[38;2;138;129;54mu[38;2;109;111;61mr[38;2;127;144;84mc[38;2;189;214;128mw[38;2;208;230;168mh[38;2;101;130;81mn[38;2;121;159;84mz[38;2;126;163;83mX[38;2;123;158;82mz[38;2;154;196;96mL[38;2;168;212;101mO[38;2;165;208;101m0[38;2;124;152;72mc[38;2;125;121;59mn[38;2;195;175;85mQ[38;2;201;173;71mL[38;2;160;122;48mv[38;2;153;119;45mn[38;2;227;206;86mm[38;2;222;209;94mw[38;2;151;140;62mc[38;2;219;208;115mq[38;2;212;201;77mO[38;2;202;189;89mO[38;2;145;133;68mc[38;2;194;185;123mZ[38;2;194;188;135mm[38;2;93;84;54m1[38;2;33;28;27m;[38;2;0;0;0m                                                                                    [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;7;6;5m.[38;2;92;91;59mt[38;2;135;131;74mv[38;2;116;105;53mj[38;2;137;123;67mu[38;2;142;128;60mv[38;2;137;124;58mu[38;2;130;116;52mx[38;2;154;138;62mc[38;2;198;182;82mQ[38;2;210;195;82mO[38;2;208;193;82mO[38;2;196;181;78mQ[38;2;193;178;84mQ[38;2;195;179;89mQ[38;2;198;183;92m0[38;2;211;196;101mZ[38;2;230;218;108mp[38;2;227;217;103mq[38;2;200;190;82m0[38;2;217;206;101mw[38;2;237;226;122mb[38;2;223;215;114mp[38;2;164;150;72mY[38;2;144;134;60mv[38;2;206;197;134mq[38;2;170;155;72mY[38;2;230;213;100mq[38;2;118;105;45mj[38;2;97;84;42m1[38;2;154;134;66mc[38;2;171;147;73mY[38;2;134;122;57mn[38;2;121;124;56mx[38;2;136;149;68mc[38;2;122;142;63mu[38;2;106;129;59mx[38;2;104;132;59mx[38;2;149;177;92mJ[38;2;194;222;147mp[38;2;112;149;83mv[38;2;116;162;80mz[38;2;124;173;77mX[38;2;136;187;83mU[38;2;144;193;91mC[38;2;154;203;96mQ[38;2;161;209;101m0[38;2;145;180;100mJ[38;2;75;82;46m-[38;2;128;120;68mn[38;2;120;98;45mj[38;2;119;84;43mt[38;2;90;60;28m+[38;2;177;165;72mJ[38;2;244;236;100mb[38;2;168;158;62mY[38;2;212;203;109mw[38;2;212;201;88mZ[38;2;178;161;82mJ[38;2;136;116;59mn[38;2;197;182;94m0[38;2;219;206;142md[38;2;158;154;125mC[38;2;14;15;12m'[38;2;0;0;0m     [38;2;11;11;11m'[38;2;46;46;46mi[38;2;64;64;64m-[38;2;66;66;66m-[38;2;65;65;65m---------------[38;2;66;66;66m-[38;2;64;64;64m-[38;2;48;48;48mi[38;2;12;12;12m'[38;2;0;0;0m  [38;2;18;18;18m^[38;2;52;52;52m~[38;2;65;65;65m-[38;2;66;66;66m-[38;2;65;65;65m---[38;2;66;66;66m-[38;2;63;63;63m_[38;2;41;41;41ml[38;2;6;6;6m.[38;2;0;0;0m       [38;2;8;8;8m.[38;2;44;44;44m![38;2;64;64;64m-[38;2;66;66;66m-[38;2;65;65;65m---[38;2;66;66;66m-[38;2;65;65;65m-[38;2;50;50;50mi[38;2;16;16;16m^[38;2;20;20;20m\"[38;2;54;54;54m~[38;2;65;65;65m-[38;2;66;66;66m-[38;2;65;65;65m---[38;2;66;66;66m-[38;2;62;62;62m_[38;2;39;39;39ml[38;2;4;4;4m [38;2;0;0;0m              [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;4;2;2m [38;2;103;102;57mj[38;2;176;175;90mL[38;2;113;99;56mj[38;2;130;116;59mn[38;2;208;200;86mO[38;2;211;204;87mZ[38;2;208;200;92mZ[38;2;192;183;88mQ[38;2;185;175;86mL[38;2;190;181;86mQ[38;2;176;165;82mJ[38;2;166;152;82mU[38;2;167;151;82mU[38;2;169;155;77mU[38;2;172;158;76mU[38;2;183;171;85mC[38;2;191;179;84mQ[38;2;203;192;91mO[38;2;208;199;92mZ[38;2;184;177;80mL[38;2;143;136;65mv[38;2;119;112;65mx[38;2;142;131;69mv[38;2;171;164;73mU[38;2;185;178;106m0[38;2;178;164;74mJ[38;2;225;208;90mw[38;2;144;141;60mc[38;2;150;170;81mU[38;2;143;172;71mY[38;2;133;159;67mz[38;2;138;174;73mY[38;2;124;165;55mv[38;2;128;165;59mc[38;2;122;156;58mv[38;2;111;142;55mn[38;2;97;121;49mj[38;2;80;97;46m1[38;2;129;151;93mX[38;2;164;196;119m0[38;2;162;200;121mO[38;2;125;166;89mX[38;2;111;152;73mv[38;2;137;178;91mU[38;2;135;171;94mU[38;2;115;147;85mc[38;2;92;121;65mr[38;2;66;88;47m-[38;2;68;85;43m-[38;2;116;132;60mn[38;2;151;161;83mY[38;2;69;64;32m+[38;2;172;169;76mJ[38;2;226;216;91mw[38;2;186;171;57mJ[38;2;221;208;89mm[38;2;215;207;82mZ[38;2;151;136;67mc[38;2;127;109;49mr[38;2;182;165;69mJ[38;2;197;182;87mQ[38;2;162;159;104mJ[38;2;22;23;17m\"[38;2;0;0;0m   [38;2;5;5;5m.[38;2;114;114;114mv[38;2;216;216;216m*[38;2;251;251;251m@[38;2;255;255;255m$$$$$$$$$$$$$$$$$$$[38;2;252;251;251m@[38;2;219;219;219m*[38;2;124;124;124mX[38;2;139;139;139mJ[38;2;227;227;227mM[38;2;253;253;253m$[38;2;255;255;255m$$$$$$$[38;2;247;248;247m@[38;2;206;206;206ma[38;2;92;92;92mr[38;2;0;0;0m    [38;2;2;2;2m [38;2;103;103;103mn[38;2;211;211;211mo[38;2;249;249;249m@[38;2;255;255;255m$$$$$$$[38;2;253;252;253m$[38;2;225;225;225mM[38;2;230;230;230mW[38;2;254;254;254m$[38;2;255;255;255m$$$$$$$[38;2;246;246;246mB[38;2;201;201;201mk[38;2;83;83;83mf[38;2;0;0;0m             [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;0;0;1m [38;2;5;5;5m.[38;2;67;67;40m+[38;2;173;171;86mC[38;2;143;129;67mv[38;2;129;113;61mn[38;2;198;188;102mO[38;2;177;166;95mC[38;2;166;154;92mU[38;2;162;150;80mY[38;2;173;161;85mJ[38;2;183;170;96mL[38;2;183;169;90mL[38;2;183;169;86mC[38;2;182;169;84mC[38;2;173;166;72mU[38;2;161;158;69mY[38;2;154;152;74mX[38;2;155;156;80mY[38;2;117;122;48mr[38;2;119;132;55mn[38;2;134;153;67mc[38;2;143;166;71mX[38;2;149;174;75mY[38;2;120;132;51mn[38;2;186;189;93m0[38;2;167;164;70mU[38;2;185;173;86mL[38;2;183;167;59mU[38;2;219;207;95mm[38;2;166;162;72mU[38;2;124;137;55mn[38;2;140;164;70mX[38;2;130;160;62mc[38;2;122;150;64mv[38;2;140;157;90mY[38;2;151;158;109mJ[38;2;170;169;131m0[38;2;191;184;144mm[38;2;192;182;142mm[38;2;189;183;146mm[38;2;187;190;148mw[38;2;148;161;109mJ[38;2;142;164;106mU[38;2;104;127;76mn[38;2;70;88;55m?[38;2;22;29;19m,[38;2;19;22;11m^[38;2;115;127;71mn[38;2;146;167;82mY[38;2;113;140;65mu[38;2;106;135;59mx[38;2;163;188;99mL[38;2;94;99;46mt[38;2;206;204;94mZ[38;2;197;187;64mL[38;2;215;200;71mO[38;2;225;206;80mm[38;2;210;191;86mO[38;2;123;101;42mj[38;2;192;176;90mQ[38;2;178;164;72mJ[38;2;168;152;70mY[38;2;145;138;76mz[38;2;20;19;16m^[38;2;0;0;0m   [38;2;111;111;111mv[38;2;255;255;255m$$$[38;2;255;253;254m$[38;2;254;248;247m@@[38;2;253;248;247m@[38;2;253;247;247m@[38;2;253;248;247m@[38;2;253;247;247m@[38;2;253;248;247m@[38;2;254;248;247m@@@@@@@@[38;2;253;247;247m@[38;2;253;247;246m@[38;2;254;252;252m$[38;2;255;255;255m$$$$$[38;2;254;255;255m$[38;2;252;253;253m$[38;2;254;247;247m@@[38;2;253;247;247m@@[38;2;252;247;248m@[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;254;254;254m$[38;2;97;97;97mx[38;2;0;0;0m   [38;2;90;90;90mj[38;2;255;255;255m$$$[38;2;253;253;252m$[38;2;254;247;247m@@@[38;2;253;247;247m@[38;2;253;247;246m@[38;2;253;251;252m$[38;2;255;255;255m$$$$[38;2;254;250;250m@[38;2;252;247;246m@[38;2;253;247;247m@@[38;2;254;247;247m@[38;2;253;248;247m@[38;2;255;255;255m$$$[38;2;251;251;251m@[38;2;61;61;61m_[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;2;2;2m [38;2;77;77;54m?[38;2;149;141;86mX[38;2;196;187;104mO[38;2;194;182;101m0[38;2;146;131;68mc[38;2;127;113;61mx[38;2;122;106;62mx[38;2;125;109;54mx[38;2;151;138;60mc[38;2;170;164;70mU[38;2;173;171;77mJ[38;2;179;184;84mL[38;2;176;188;82mL[38;2;164;182;75mJ[38;2;156;181;68mU[38;2;154;184;71mU[38;2;146;176;69mY[38;2;157;190;75mJ[38;2;174;211;84m0[38;2;173;214;81m0[38;2;169;212;75mQ[38;2;167;210;69mL[38;2;163;205;68mC[38;2;153;191;69mU[38;2;148;175;67mY[38;2;141;146;69mc[38;2;138;129;63mv[38;2;149;133;63mc[38;2;180;158;63mU[38;2;228;208;86mw[38;2;235;221;89mq[38;2;224;215;92mw[38;2;188;182;80mL[38;2;179;171;91mL[38;2;194;178;131mZ[38;2;252;234;194mM[38;2;255;241;197mW[38;2;255;242;200mW[38;2;200;181;144mw[38;2;205;190;158mp[38;2;255;248;215m8[38;2;238;223;193m*[38;2;144;138;109mY[38;2;104;104;80mx[38;2;16;16;13m^[38;2;16;9;7m'[38;2;167;130;100mY[38;2;237;184;119mq[38;2;213;174;101mO[38;2;164;148;78mY[38;2;147;164;76mY[38;2;141;162;77mX[38;2;149;152;71mX[38;2;211;203;84mZ[38;2;212;200;73mO[38;2;220;204;83mZ[38;2;175;153;74mU[38;2;139;117;51mn[38;2;166;150;72mY[38;2;138;124;56mu[38;2;170;154;80mU[38;2;173;154;76mU[38;2;146;138;86mz[38;2;8;8;8m.[38;2;0;0;0m [38;2;0;0;1m [38;2;0;0;0m [38;2;161;161;161mO[38;2;255;255;255m$$[38;2;250;255;255m$[38;2;225;169;173md[38;2;248;44;51mv[38;2;253;45;52mc[38;2;253;45;53mc[38;2;252;45;52mc[38;2;252;44;53mccc[38;2;253;43;53mc[38;2;253;43;52mccc[38;2;252;41;52mc[38;2;252;40;53mc[38;2;252;40;52mvv[38;2;252;40;51mv[38;2;250;38;46mv[38;2;224;151;155mw[38;2;248;254;254m$[38;2;255;255;255m$$$$[38;2;235;233;233mW[38;2;236;82;91mU[38;2;250;38;47mv[38;2;250;39;51mv[38;2;248;39;50mv[38;2;247;38;50mv[38;2;246;39;46mv[38;2;228;143;148mm[38;2;246;254;254m@[38;2;255;255;255m$$[38;2;234;234;234m&[38;2;38;38;38ml[38;2;0;0;0m  [38;2;146;146;146mC[38;2;255;255;255m$$[38;2;251;255;255m$[38;2;218;177;178md[38;2;232;39;49mu[38;2;239;38;48mu[38;2;238;39;49muu[38;2;236;37;43mn[38;2;219;134;139mO[38;2;247;252;253m@[38;2;255;255;255m$$[38;2;242;248;248mB[38;2;216;112;117mL[38;2;234;37;41mn[38;2;233;39;49mu[38;2;232;38;47mn[38;2;233;38;46mn[38;2;223;48;55mu[38;2;222;201;202ma[38;2;254;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;56;50;30m![38;2;190;171;94mQ[38;2;192;173;79mL[38;2;166;148;61mX[38;2;159;138;56mc[38;2;143;128;49mu[38;2;112;106;40mf[38;2;130;143;57mv[38;2;180;212;88mO[38;2;191;228;91mm[38;2;173;209;78mQ[38;2;154;186;75mJ[38;2;151;180;74mU[38;2;159;190;78mC[38;2;178;216;81m0[38;2;183;228;83mO[38;2;157;197;74mC[38;2;121;154;55mv[38;2;113;141;52mn[38;2;116;141;57mn[38;2;119;139;60mu[38;2;121;134;62mn[38;2;129;138;70mv[38;2;126;135;67mu[38;2;127;133;77mv[38;2;129;124;86mv[38;2;142;129;97mz[38;2;167;151;105mJ[38;2;156;139;77mX[38;2;157;139;71mz[38;2;163;148;68mX[38;2;201;189;81m0[38;2;247;235;92md[38;2;255;243;98mk[38;2;171;153;77mU[38;2;221;202;165mb[38;2;255;237;199mW[38;2;249;230;187m#[38;2;165;147;108mJ[38;2;163;145;112mJ[38;2;228;208;171mh[38;2;213;191;149mp[38;2;176;156;117mL[38;2;149;132;101mX[38;2;112;101;83mx[38;2;33;19;15m\"[38;2;152;116;85mc[38;2;188;142;84mJ[38;2;163;126;70mz[38;2;135;102;63mx[38;2;91;70;42m-[38;2;137;127;63mu[38;2;188;172;78mC[38;2;176;165;58mU[38;2;183;184;73mC[38;2;153;157;65mX[38;2;95;91;42m1[38;2;125;115;63mn[38;2;94;80;38m?[38;2;93;77;44m?[38;2;173;155;74mU[38;2;221;200;99mm[38;2;132;126;73mv[38;2;6;7;7m.[38;2;2;2;3m [38;2;0;0;0m  [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;255;254m$[38;2;209;141;144mO[38;2;250;0;9mf[38;2;255;2;12mj[38;2;255;3;12mj[38;2;254;2;11mj[38;2;254;2;13mj[38;2;255;0;11mj[38;2;253;0;7mf[38;2;254;0;6mf[38;2;254;0;5mfff[38;2;253;0;5mf[38;2;253;0;4mffff[38;2;250;0;0mf[38;2;206;114;119mC[38;2;244;252;252m@[38;2;255;255;255m$$$[38;2;245;252;252m@[38;2;219;119;125mQ[38;2;247;0;6mf[38;2;252;0;10mj[38;2;251;0;10mj[38;2;249;0;10mf[38;2;248;0;9mf[38;2;249;0;6mf[38;2;234;16;27mr[38;2;221;191;193mk[38;2;254;255;255m$[38;2;255;255;255m$$[38;2;185;185;185mp[38;2;5;5;5m.[38;2;0;0;0m [38;2;157;157;157m0[38;2;255;255;255m$$[38;2;249;255;254m$[38;2;199;149;151mZ[38;2;231;0;6mt[38;2;240;0;7mt[38;2;238;0;8mtt[38;2;236;0;1mt[38;2;202;100;105mU[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;233;241;240m8[38;2;198;73;79mc[38;2;233;0;0m1[38;2;232;0;8mt[38;2;231;0;6mt[38;2;231;0;4mt[38;2;216;4;13m1[38;2;203;177;180mp[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;33;29;22m;[38;2;136;120;71mu[38;2;145;126;60mv[38;2;135;120;52mn[38;2;139;130;57mu[38;2;133;133;59mu[38;2;144;160;70mX[38;2;184;219;90mO[38;2;142;179;69mY[38;2;97;126;50mj[38;2;127;156;67mc[38;2;187;220;93mZ[38;2;198;235;91mw[38;2;186;225;80mO[38;2;163;196;75mC[38;2;122;146;59mu[38;2;85;94;46m1[38;2;75;75;58m?[38;2;86;84;72mt[38;2;41;38;35ml[38;2;26;22;20m\"[38;2;23;18;17m\"[38;2;30;23;23m,[38;2;37;32;27mI[38;2;46;42;33ml[38;2;60;54;43m~[38;2;71;63;51m_[38;2;79;70;57m-[38;2;85;76;60m?[38;2;120;110;80mn[38;2;128;117;88mv[38;2;96;83;53m1[38;2;164;145;72mX[38;2;235;220;88mq[38;2;211;198;89mZ[38;2;180;163;108mL[38;2;251;231;185m#[38;2;188;163;120m0[38;2;139;114;73mu[38;2;109;85;48mt[38;2;131;105;75mn[38;2;184;161;127m0[38;2;210;187;151mq[38;2;174;154;112mC[38;2;176;159;118mQ[38;2;126;110;86mu[38;2;37;20;16m,[38;2;59;44;31m![38;2;81;64;42m_[38;2;100;81;41m1[38;2;173;150;83mU[38;2;170;136;70mX[38;2;194;153;88mC[38;2;178;153;80mU[38;2;143;140;69mc[38;2;138;152;83mX[38;2;51;61;32mi[38;2;51;47;32m![38;2;79;66;40m_[38;2;157;139;72mz[38;2;193;176;69mC[38;2;223;208;106mq[38;2;142;130;60mv[38;2;182;181;95mQ[38;2;110;112;70mx[38;2;2;1;1m [38;2;0;0;0m [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;254;5;14mj[38;2;197;51;58mn[38;2;185;108;112mU[38;2;192;111;115mJ[38;2;192;110;115mJ[38;2;192;111;115mJ[38;2;191;110;114mJ[38;2;192;109;114mJJJJ[38;2;192;109;113mJ[38;2;196;114;118mC[38;2;217;189;189mk[38;2;251;254;253m$[38;2;255;255;255m$$[38;2;252;255;255m$[38;2;221;181;183mb[38;2;238;13;24mj[38;2;252;0;14mj[38;2;251;0;15mjj[38;2;251;0;14mj[38;2;248;1;14mjj[38;2;248;0;7mf[38;2;224;58;69mc[38;2;234;232;234mW[38;2;255;255;255m$$$[38;2;117;117;117mc[38;2;0;0;0m [38;2;156;156;156m0[38;2;255;255;255m$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;20;20;17m\"[38;2;116;118;72mn[38;2;160;163;84mU[38;2;174;186;90mL[38;2;173;198;89mQ[38;2;158;186;80mJ[38;2;118;142;67mu[38;2;70;90;35m-[38;2;93;115;51mf[38;2;155;188;79mJ[38;2;188;228;89mZ[38;2;166;202;73mL[38;2;124;151;60mv[38;2;106;125;59mx[38;2;98;103;67mj[38;2;82;74;47m-[38;2;122;103;61mr[38;2;120;92;57mj[38;2;155;130;107mY[38;2;183;166;144mO[38;2;185;175;149mZ[38;2;164;156;130mL[38;2;146;136;114mY[38;2;139;132;112mX[38;2;144;136;117mY[38;2;158;151;132mL[38;2;177;169;149mZ[38;2;136;128;110mX[38;2;73;67;56m-[38;2;24;20;17m\"[38;2;11;8;9m.[38;2;7;2;3m [38;2;85;76;50m?[38;2;173;162;80mJ[38;2;209;194;85mO[38;2;201;186;88m0[38;2;185;163;99mL[38;2;142;116;68mu[38;2;144;110;64mu[38;2;154;114;60mu[38;2;198;161;110m0[38;2;149;128;100mX[38;2;224;215;192ma[38;2;183;168;130mO[38;2;178;156;116mL[38;2;221;206;164mk[38;2;55;45;35m![38;2;63;48;32mi[38;2;128;99;61mx[38;2;163;126;66mc[38;2;185;139;74mY[38;2;211;164;100m0[38;2;243;197;120mp[38;2;173;141;88mU[38;2;64;50;30mi[38;2;17;13;10m'[38;2;0;0;0m [38;2;28;24;12m\"[38;2;155;143;74mX[38;2;192;176;73mL[38;2;200;194;97mO[38;2;129;123;69mu[38;2;141;131;64mv[38;2;209;202;97mZ[38;2;131;128;81mv[38;2;2;1;2m [38;2;0;0;0m [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;253;0;10mj[38;2;205;116;119mC[38;2;235;252;252mB[38;2;249;255;255m$$$$$$$$$$[38;2;254;255;255m$[38;2;255;255;255m$$$[38;2;231;228;227mM[38;2;229;51;60mv[38;2;252;0;8mf[38;2;251;1;15mj[38;2;251;0;15mj[38;2;247;0;13mf[38;2;227;1;13mt[38;2;250;0;12mj[38;2;247;1;16mj[38;2;248;0;16mj[38;2;246;0;10mf[38;2;218;118;125mQ[38;2;244;252;252m@[38;2;255;255;255m$$[38;2;242;242;242m8[38;2;42;42;42m![38;2;149;149;149mL[38;2;255;255;255m$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                        [38;2;1;1;2m [38;2;44;51;28ml[38;2;130;149;81mz[38;2;165;194;86mL[38;2;170;200;86mQ[38;2;146;174;73mY[38;2;109;137;62mn[38;2;77;99;44m?[38;2;92;115;47mf[38;2;156;189;76mJ[38;2;183;223;86mO[38;2;158;198;74mC[38;2;109;138;52mx[38;2;100;105;53mf[38;2;114;109;58mr[38;2;128;122;64mn[38;2;83;69;39m_[38;2;175;156;117mL[38;2;231;203;145mb[38;2;190;156;100mL[38;2;138;107;60mn[38;2;115;89;51mf[38;2;117;98;70mr[38;2;151;138;114mU[38;2;172;159;135mQ[38;2;182;172;147mZ[38;2;187;177;152mm[38;2;196;186;161mq[38;2;204;193;168md[38;2;218;205;172mk[38;2;210;197;163md[38;2;176;164;136m0[38;2;143;130;112mY[38;2;115;103;89mn[38;2;65;54;45m~[38;2;110;95;60mj[38;2;154;132;78mz[38;2;155;138;72mz[38;2;185;176;93mQ[38;2;122;108;67mx[38;2;57;37;25ml[38;2;139;108;64mn[38;2;195;158;96mL[38;2;132;108;69mn[38;2;196;187;161mq[38;2;201;185;158mq[38;2;132;118;97mc[38;2;87;82;69mt[38;2;5;2;1m [38;2;95;79;61mt[38;2;154;127;95mX[38;2;100;68;41m?[38;2;135;101;68mn[38;2;130;106;75mn[38;2;61;49;31mi[38;2;15;7;7m.[38;2;16;11;10m'[38;2;18;14;15m^[38;2;32;27;22m,[38;2;94;87;45m1[38;2;176;167;81mJ[38;2;170;164;76mU[38;2;123;122;72mn[38;2;144;140;96mX[38;2;159;146;72mX[38;2;183;171;98mL[38;2;119;114;88mu[38;2;0;0;0m  [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;253;0;10mj[38;2;210;116;119mL[38;2;243;253;253m@[38;2;255;255;255m$$$$$$$$$$$$$[38;2;243;250;251m@[38;2;220;110;118mL[38;2;249;0;8mf[38;2;253;0;15mj[38;2;251;0;15mj[38;2;252;0;11mj[38;2;210;34;44mx[38;2;154;94;97mc[38;2;239;6;20mj[38;2;249;0;14mj[38;2;248;0;16mj[38;2;249;0;13mj[38;2;236;13;24mj[38;2;221;181;184mb[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;186;186;186mp[38;2;164;164;164mO[38;2;255;255;255m$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                      [38;2;0;0;1m [38;2;0;0;0m [38;2;32;38;24m;[38;2;153;176;102mC[38;2;151;183;80mJ[38;2;121;156;58mv[38;2;111;144;60mn[38;2;113;143;63mu[38;2;139;172;70mX[38;2;181;219;84mO[38;2;188;228;87mZ[38;2;149;185;69mU[38;2;105;132;49mr[38;2;61;68;33m~[38;2;94;88;53mt[38;2;152;136;64mc[38;2;182;173;86mL[38;2;173;161;89mJ[38;2;113;92;53mf[38;2;210;187;137mw[38;2;255;227;168m*[38;2;248;218;160ma[38;2;213;184;128mw[38;2;163;132;82mX[38;2;115;90;60mj[38;2;78;63;52m-[38;2;70;61;58m_[38;2;78;72;70m?[38;2;100;97;93mx[38;2;105;101;97mn[38;2;109;106;99mn[38;2;123;119;111mc[38;2;108;103;97mn[38;2;97;90;83mj[38;2;94;87;80mj[38;2;113;107;98mu[38;2;109;101;92mx[38;2;89;80;68mt[38;2;72;62;52m_[38;2;107;95;58mf[38;2;159;143;80mX[38;2;136;125;79mv[38;2;5;0;0m [38;2;21;11;9m'[38;2;79;59;39m+[38;2;92;71;49m?[38;2;145;131;110mY[38;2;127;113;96mv[38;2;28;23;17m\"[38;2;0;0;0m [38;2;2;0;3m [38;2;10;3;1m [38;2;47;37;30ml[38;2;60;47;42mi[38;2;70;56;46m+[38;2;94;80;66mt[38;2;126;111;90mu[38;2;178;160;129mQ[38;2;205;187;152mq[38;2;127;111;85mu[38;2;109;97;62mj[38;2;139;128;65mv[38;2;134;121;52mn[38;2;192;182;119mO[38;2;146;145;113mU[38;2;130;132;111mX[38;2;99;96;58mf[38;2;66;61;41m+[38;2;14;14;11m'[38;2;0;0;0m  [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;252;1;12mj[38;2;208;110;114mC[38;2;238;238;239m8[38;2;250;243;244mB[38;2;250;243;243mB[38;2;249;243;243mBBBBBB[38;2;250;245;246m@[38;2;254;253;254m$[38;2;253;254;254m$[38;2;254;255;255m$[38;2;251;255;255m$[38;2;220;173;176md[38;2;241;9;22mj[38;2;253;0;12mj[38;2;252;0;15mj[38;2;253;0;14mj[38;2;241;3;14mf[38;2;193;139;144m0[38;2;210;224;223m*[38;2;202;72;78mc[38;2;249;0;9mf[38;2;248;0;16mjj[38;2;249;0;9mf[38;2;224;50;59mv[38;2;230;227;228mM[38;2;255;255;255m$$$[38;2;241;241;241m8[38;2;255;255;255m$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                        [38;2;12;14;10m'[38;2;77;92;53m1[38;2;125;150;68mv[38;2;154;185;77mJ[38;2;173;206;92m0[38;2;181;215;90mO[38;2;183;217;82mO[38;2;161;196;73mC[38;2;107;137;51mx[38;2;62;78;37m+[38;2;57;63;30mi[38;2;120;111;52mr[38;2;179;164;75mJ[38;2;179;168;78mJ[38;2;149;134;57mv[38;2;114;91;35mt[38;2;153;127;87mz[38;2;241;217;162ma[38;2;253;223;167mo[38;2;254;221;166mo[38;2;246;216;161ma[38;2;212;182;128mw[38;2;147;119;80mc[38;2;108;84;62mf[38;2;54;36;22ml[38;2;45;36;30ml[38;2;104;102;100mn[38;2;144;143;145mC[38;2;106;104;106mn[38;2;103;101;98mx[38;2;72;71;65m?[38;2;63;63;56m_[38;2;84;86;80mf[38;2;139;140;136mJ[38;2;135;130;134mU[38;2;84;81;84mf[38;2;66;64;65m-[38;2;77;64;42m_[38;2;186;164;89mC[38;2;101;83;47m1[38;2;17;11;8m'[38;2;49;47;37m![38;2;68;58;45m+[38;2;140;122;102mz[38;2;184;165;135mO[38;2;140;126;106mX[38;2;17;16;12m^[38;2;0;0;0m [38;2;11;11;8m'[38;2;113;111;104mu[38;2;159;156;147mQ[38;2;184;179;169mw[38;2;190;180;167mq[38;2;193;182;165mq[38;2;174;163;145mO[38;2;121;111;94mu[38;2;74;65;46m_[38;2;121;112;76mn[38;2;121;112;71mn[38;2;111;98;50mf[38;2;141;128;55mu[38;2;209;203;120mw[38;2;174;178;135mO[38;2;77;84;81mt[38;2;2;4;5m [38;2;0;0;0m    [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;254;7;16mr[38;2;253;6;16mj[38;2;244;22;31mx[38;2;246;42;50mv[38;2;249;41;51mvv[38;2;249;40;51mvvv[38;2;248;39;51mv[38;2;248;38;50mv[38;2;249;36;48mv[38;2;241;50;61mc[38;2;230;203;206mo[38;2;252;255;255m$[38;2;255;255;255m$[38;2;228;223;222mM[38;2;231;45;55mv[38;2;254;0;10mj[38;2;252;0;15mjj[38;2;254;0;8mj[38;2;203;66;73mv[38;2;221;228;227mM[38;2;252;255;255m$[38;2;200;180;183mp[38;2;225;18;28mj[38;2;249;0;14mj[38;2;248;0;16mj[38;2;248;0;15mj[38;2;246;0;8mf[38;2;218;108;114mC[38;2;242;250;250m@[38;2;255;255;255m$$$$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                        [38;2;0;0;1m [38;2;48;55;35mi[38;2;140;159;95mY[38;2;197;214;143mp[38;2;213;224;175mh[38;2;206;214;176mk[38;2;181;183;143mZ[38;2;166;169;125mQ[38;2;133;132;98mz[38;2;96;89;52mt[38;2;176;170;86mC[38;2;198;181;78mQ[38;2;163;143;51mz[38;2;155;137;53mc[38;2;179;156;68mU[38;2;195;166;87mL[38;2;133;106;58mx[38;2;220;193;149mp[38;2;232;203;156mk[38;2;218;191;147mp[38;2;205;180;137mw[38;2;191;168;128mO[38;2;171;146;109mC[38;2;153;125;90mz[38;2;136;105;70mn[38;2;122;90;54mj[38;2;130;104;67mx[38;2;134;116;91mv[38;2;117;106;95mu[38;2;108;102;99mn[38;2;113;110;106mu[38;2;131;128;123mX[38;2;155;154;146mQ[38;2;160;160;153m0[38;2;149;148;139mC[38;2;92;90;88mj[38;2;39;38;39ml[38;2;78;64;33m+[38;2;201;178;98m0[38;2;120;94;59mj[38;2;191;176;147mm[38;2;238;230;202m#[38;2;208;196;170md[38;2;194;175;137mZ[38;2;255;238;190mM[38;2;224;207;174mk[38;2;33;29;23m;[38;2;12;12;12m'[38;2;93;94;90mr[38;2;116;115;112mv[38;2;107;106;103mn[38;2;82;82;79mt[38;2;69;70;67m-[38;2;72;73;70m?[38;2;37;37;34mI[38;2;35;35;32mI[38;2;64;61;58m_[38;2;82;73;71m1[38;2;64;53;29mi[38;2;136;126;66mu[38;2;141;135;61mv[38;2;166;166;109mL[38;2;91;97;74mj[38;2;16;18;16m^[38;2;0;0;0m     [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;254;7;16mr[38;2;254;7;17mr[38;2;255;2;12mj[38;2;255;0;7mj[38;2;255;0;8mj[38;2;255;0;7mjjj[38;2;255;0;8mj[38;2;255;0;7mj[38;2;255;0;6mj[38;2;255;0;3mf[38;2;244;0;12mf[38;2;212;177;180md[38;2;253;255;255m$[38;2;242;249;248mB[38;2;220;102;110mC[38;2;251;0;9mf[38;2;253;0;16mj[38;2;252;0;15mj[38;2;255;0;12mj[38;2;228;18;30mr[38;2;200;180;181mp[38;2;251;255;255m$[38;2;255;255;255m$[38;2;237;248;248mB[38;2;192;117;121mC[38;2;242;1;12mf[38;2;249;0;16mj[38;2;248;0;16mj[38;2;249;0;14mj[38;2;235;9;20mj[38;2;219;172;174md[38;2;251;255;255m$[38;2;255;255;255m$$$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;113;113;113mv[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;44;46;44m![38;2;194;199;184mb[38;2;249;247;226m8[38;2;246;240;220m&[38;2;239;233;213mM[38;2;251;245;224m8[38;2;214;209;186mh[38;2;214;205;176mk[38;2;226;213;173mh[38;2;129;112;76mn[38;2;134;121;59mn[38;2;191;181;75mL[38;2;197;179;74mL[38;2;159;134;57mc[38;2;126;104;46mr[38;2;95;76;56m1[38;2;211;198;183mk[38;2;240;230;214mM[38;2;230;225;210m#[38;2;232;227;213mM[38;2;228;224;212m#[38;2;213;206;191mh[38;2;208;196;177mb[38;2;163;137;109mU[38;2;138;99;54mx[38;2;151;108;53mn[38;2;178;144;94mJ[38;2;189;170;134mO[38;2;205;190;174md[38;2;216;207;192mh[38;2;178;171;156mZ[38;2;153;146;132mC[38;2;115;105;93mn[38;2;69;58;50m+[38;2;38;33;28mI[38;2;28;23;10m\"[38;2;107;83;41m1[38;2;181;152;84mJ[38;2;214;192;152mp[38;2;254;243;213m&[38;2;255;249;237m@@[38;2;191;178;147mm[38;2;218;198;151md[38;2;199;181;139mm[38;2;91;82;66mt[38;2;27;23;21m,[38;2;76;74;73m1[38;2;82;82;79mt[38;2;69;69;66m-[38;2;49;51;47mi[38;2;72;74;70m?[38;2;96;97;94mr[38;2;82;81;78mt[38;2;185;183;180mq[38;2;163;159;154m0[38;2;40;34;27mI[38;2;138;127;72mv[38;2;126;107;60mx[38;2;77;71;52m-[38;2;25;26;22m,[38;2;0;0;0m       [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;254;7;16mr[38;2;254;6;16mr[38;2;214;28;37mr[38;2;200;56;62mu[38;2;206;57;65mu[38;2;205;57;65muu[38;2;205;56;64muu[38;2;205;55;63muu[38;2;205;54;62mu[38;2;207;71;79mz[38;2;221;203;204ma[38;2;249;255;255m$[38;2;221;166;169mp[38;2;242;7;20mj[38;2;254;0;13mj[38;2;253;1;16mj[38;2;251;0;15mj[38;2;247;1;12mf[38;2;195;92;99mY[38;2;226;224;225mM[38;2;247;237;238m8[38;2;246;236;237m8[38;2;247;238;238m8[38;2;205;197;196mk[38;2;209;41;52mx[38;2;250;0;12mj[38;2;248;0;16mjj[38;2;247;0;8mf[38;2;224;42;52mu[38;2;229;221;222mM[38;2;255;255;255m$$$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;109;109;109mu[38;2;0;0;0m            [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;52;52;51m~[38;2;236;235;225mW[38;2;204;198;177mb[38;2;104;92;73mj[38;2;112;94;74mr[38;2;190;171;141mZ[38;2;247;237;201mM[38;2;221;212;181mh[38;2;221;206;171mk[38;2;227;212;183ma[38;2;104;90;65mf[38;2;111;98;45mf[38;2;179;162;81mJ[38;2;92;70;26m_[38;2;141;120;77mv[38;2;171;159;129mQ[38;2;148;146;131mJ[38;2;250;249;243m@[38;2;255;253;247m@[38;2;255;252;248m@[38;2;254;253;247m@[38;2;255;255;243m@[38;2;231;222;197m*[38;2;202;173;120mZ[38;2;206;158;88mL[38;2;198;145;71mJ[38;2;198;146;77mJ[38;2;193;147;85mJ[38;2;177;136;88mU[38;2;172;140;95mU[38;2;138;111;71mu[38;2;91;68;35m-[38;2;85;64;37m_[38;2;72;51;36m~[38;2;66;47;25mi[38;2;142;124;64mv[38;2;201;173;91mQ[38;2;192;169;112m0[38;2;249;241;215m&[38;2;255;252;241m@[38;2;254;250;241m@[38;2;255;251;240m@[38;2;249;241;216m&[38;2;190;171;130mO[38;2;153;131;92mX[38;2;140;126;101mz[38;2;88;79;65m1[38;2;50;44;40m![38;2;3;2;1m [38;2;51;50;48mi[38;2;116;111;101mu[38;2;165;154;135mQ[38;2;188;176;154mm[38;2;212;205;190mh[38;2;255;255;248m$[38;2;171;169;161mZ[38;2;89;82;48m?[38;2;144;128;79mc[38;2;80;65;47m-[38;2;19;17;19m^[38;2;0;0;0m        [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;253;1;11mj[38;2;198;108;111mJ[38;2;219;235;235mW[38;2;232;240;240m&[38;2;231;240;240m&[38;2;232;240;240m&[38;2;233;241;241m88[38;2;232;240;240m&[38;2;231;240;240m&&[38;2;237;245;245m8[38;2;250;255;254m$[38;2;228;217;218m#[38;2;231;40;50mu[38;2;254;0;10mj[38;2;253;1;16mjj[38;2;252;0;15mj[38;2;248;2;15mj[38;2;236;21;32mx[38;2;242;30;42mn[38;2;243;29;42mn[38;2;241;29;41mnn[38;2;238;29;40mn[38;2;236;13;25mj[38;2;249;1;14mj[38;2;248;0;16mjj[38;2;246;1;13mf[38;2;245;0;8mf[38;2;218;97;104mJ[38;2;241;248;246mB[38;2;255;255;255m$$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;179;181md[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;146;146;146mC[38;2;58;58;58m+[38;2;59;59;59m++++++[38;2;52;52;52m~[38;2;25;25;25m,[38;2;0;0;0m   [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;46;46;45m![38;2;220;220;211m*[38;2;88;79;69mt[38;2;144;123;83mc[38;2;223;188;141mp[38;2;104;69;48m?[38;2;159;138;115mU[38;2;247;237;203mW[38;2;226;217;188ma[38;2;215;203;169mb[38;2;216;195;155md[38;2;143;122;71mv[38;2;122;103;48mj[38;2;112;96;49mf[38;2;206;185;137mw[38;2;254;237;190mM[38;2;206;195;159mp[38;2;210;203;182mk[38;2;253;248;235mB[38;2;254;249;239m@[38;2;255;251;237m@[38;2;255;251;229mB[38;2;213;201;165mb[38;2;228;200;134mp[38;2;251;200;122md[38;2;249;191;111mp[38;2;247;186;106mqq[38;2;220;163;86m0[38;2;192;141;66mU[38;2;185;138;72mY[38;2;149;108;54mn[38;2;141;103;55mx[38;2;133;97;55mr[38;2;120;87;42mf[38;2;173;143;79mY[38;2;229;199;137md[38;2;250;233;194mM[38;2;255;254;234m@[38;2;255;255;250m$[38;2;255;255;248m$[38;2;255;255;243m@[38;2;255;250;228mB[38;2;191;175;145mm[38;2;171;146;112mC[38;2;231;208;169mh[38;2;195;176;141mm[38;2;160;146;122mC[38;2;60;51;42m~[38;2;44;31;18m;[38;2;137;109;67mn[38;2;204;156;89mL[38;2;210;153;86mL[38;2;237;209;155mk[38;2;255;250;229mB[38;2;141;133;118mY[38;2;134;125;71mv[38;2;81;73;41m-[38;2;14;14;13m'[38;2;0;0;0m         [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;209;143;146mZ[38;2;250;5;14mj[38;2;255;7;16mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;253;0;10mj[38;2;211;116;119mL[38;2;244;252;252m@[38;2;255;255;255m$$$[38;2;254;254;254m$[38;2;251;251;251m@[38;2;254;254;254m$[38;2;255;255;255m$$$[38;2;240;247;245mB[38;2;222;94;102mJ[38;2;252;0;8mf[38;2;254;1;16mj[38;2;253;1;16mjj[38;2;255;0;12mj[38;2;255;0;9mj[38;2;255;0;6mj[38;2;255;0;5mff[38;2;253;0;4mff[38;2;253;0;5mf[38;2;253;0;9mj[38;2;252;0;11mj[38;2;250;0;15mj[38;2;248;0;16mj[38;2;246;0;13mf[38;2;247;0;11mf[38;2;237;5;16mf[38;2;218;162;164mq[38;2;250;255;255m$[38;2;255;255;255m$$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;11mt[38;2;231;0;9mt[38;2;217;9;18mt[38;2;204;181;182md[38;2;254;255;255m$[38;2;255;255;255m$$$$$$$$$$[38;2;254;254;254m$[38;2;235;235;235m&[38;2;174;174;174mw[38;2;46;46;46mi[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;41;40;42ml[38;2;226;226;222mM[38;2;146;139;125mU[38;2;163;143;100mU[38;2;243;207;151mk[38;2;148;111;70mu[38;2;159;126;89mX[38;2;160;141;117mJ[38;2;242;237;211mW[38;2;233;221;194m*[38;2;236;218;178ma[38;2;204;187;129mm[38;2;157;137;88mX[38;2;229;211;160mk[38;2;254;234;189mM[38;2;253;235;191mM[38;2;252;237;199mW[38;2;242;230;200mM[38;2;251;244;220m8[38;2;254;247;229mB[38;2;255;248;231mB[38;2;251;244;218m&[38;2;215;199;161md[38;2;246;220;161ma[38;2;254;214;143mh[38;2;254;207;132mk[38;2;252;203;123mb[38;2;247;196;114mp[38;2;245;193;109mq[38;2;241;190;103mw[38;2;228;182;101mm[38;2;188;145;77mU[38;2;175;133;68mX[38;2;176;132;73mX[38;2;148;105;58mn[38;2;138;104;59mx[38;2;199;171;124mO[38;2;231;214;170mh[38;2;248;242;213m&[38;2;222;218;201mo[38;2;188;179;161mw[38;2;157;144;124mJ[38;2;126;108;89mu[38;2;104;80;59mt[38;2;99;74;55m1[38;2;105;85;64mf[38;2;124;106;83mn[38;2;127;108;80mn[38;2;121;99;77mx[38;2;132;99;66mx[38;2;232;191;125mq[38;2;253;198;121md[38;2;249;183;105mq[38;2;234;182;109mw[38;2;209;190;152mp[38;2;109;99;78mr[38;2;114;107;78mx[38;2;24;22;16m\"[38;2;0;0;0m          [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;253;0;10mj[38;2;210;115;118mL[38;2;242;250;250m@[38;2;255;255;255m$$[38;2;213;213;213mo[38;2;45;45;45m![38;2;64;64;64m-[38;2;231;231;231mW[38;2;255;255;255m$$[38;2;251;255;255m$[38;2;220;159;162mq[38;2;245;5;17mj[38;2;254;0;14mj[38;2;253;1;16mj[38;2;252;1;17mj[38;2;253;0;14mj[38;2;210;28;39mr[38;2;199;61;69mu[38;2;204;63;70mv[38;2;203;63;70mvv[38;2;202;63;70mvv[38;2;201;63;70mv[38;2;201;63;71mv[38;2;194;56;64mn[38;2;223;13;25mj[38;2;250;0;13mj[38;2;246;0;13mff[38;2;245;0;10mf[38;2;226;35;44mn[38;2;227;215;215m*[38;2;254;255;255m$[38;2;255;255;255m$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;12mt[38;2;230;0;9mt[38;2;217;9;19mt[38;2;201;171;174mq[38;2;247;245;246mB[38;2;249;245;245mB[38;2;249;244;245mB[38;2;249;245;245mB[38;2;250;245;246m@@@@[38;2;249;245;246mBB[38;2;251;249;249m@[38;2;255;255;255m$$$[38;2;224;224;224mM[38;2;27;27;27m,[38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;9;9;11m.[38;2;143;146;145mC[38;2;229;229;222mM[38;2;129;117;90mv[38;2;228;202;154mb[38;2;152;119;75mc[38;2;213;173;110mZ[38;2;113;86;60mf[38;2;74;69;64m?[38;2;217;208;192mh[38;2;255;245;219m8[38;2;200;186;151mq[38;2;213;197;157md[38;2;254;235;187mM[38;2;252;233;186m#[38;2;254;236;200mW[38;2;253;237;206mW[38;2;254;240;213m&[38;2;253;242;218m&[38;2;254;244;221m8[38;2;255;246;222m8[38;2;247;239;211mW[38;2;223;206;165mk[38;2;251;226;172m*[38;2;253;224;161mo[38;2;253;220;152ma[38;2;252;216;149mh[38;2;250;214;146mh[38;2;249;214;141mk[38;2;249;212;134mk[38;2;249;212;137mk[38;2;240;205;141mb[38;2;205;173;111mO[38;2;191;156;93mC[38;2;163;126;67mc[38;2;167;132;73mX[38;2;164;129;67mz[38;2;183;154;97mC[38;2;158;139;102mU[38;2;80;65;49m-[38;2;75;55;42m+[38;2;79;54;34m+[38;2;85;57;32m+[38;2;114;84;54mf[38;2;95;73;48m?[38;2;53;40;27ml[38;2;44;38;26mI[38;2;94;82;75mf[38;2;83;59;43m_[38;2;210;175;126mm[38;2;254;211;144mh[38;2;250;203;131mb[38;2;251;202;131mb[38;2;237;200;131md[38;2;110;93;63mj[38;2;93;86;80mf[38;2;59;54;54m+[38;2;0;0;1m [38;2;0;0;0m          [38;2;159;159;159m0[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;143;146mZ[38;2;250;5;14mj[38;2;255;7;17mr[38;2;255;8;17mr[38;2;255;7;16mr[38;2;253;0;10mj[38;2;210;115;118mL[38;2;242;250;250m@[38;2;255;255;255m$$[38;2;202;202;202mh[38;2;0;0;0m [38;2;143;143;143mC[38;2;255;255;255m$$[38;2;254;255;255m$[38;2;227;212;213m*[38;2;234;35;46mn[38;2;254;0;12mj[38;2;253;1;16mjj[38;2;254;0;13mj[38;2;226;20;32mr[38;2;192;176;177mq[38;2;231;244;243m8[38;2;235;245;244m8[38;2;236;246;245m8[38;2;237;247;246mBB[38;2;237;246;245m8[38;2;235;245;244m8[38;2;236;245;244m8[38;2;222;237;236mW[38;2;186;122;124mC[38;2;239;1;11mf[38;2;247;0;13mf[38;2;246;0;13mf[38;2;245;0;14mf[38;2;244;0;6mf[38;2;217;87;95mU[38;2;239;245;246mB[38;2;255;255;255m$[38;2;249;255;254m$[38;2;200;151;153mZ[38;2;232;0;11mt[38;2;241;0;12mf[38;2;239;0;13mf[38;2;238;0;13mf[38;2;236;0;6mt[38;2;203;103;108mJ[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;234;241;241m8[38;2;200;77;83mz[38;2;233;0;5mt[38;2;232;0;13mt[38;2;231;0;12mt[38;2;231;0;11mt[38;2;227;2;13mt[38;2;221;27;37mr[38;2;226;39;48mn[38;2;225;39;48mn[38;2;224;39;47mnn[38;2;223;39;47mnn[38;2;222;39;47mnn[38;2;221;39;46mn[38;2;222;38;43mn[38;2;210;68;73mc[38;2;230;225;225mM[38;2;254;255;255m$[38;2;255;255;255m$$[38;2;64;64;64m-[38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;6;7;7m.[38;2;126;128;126mX[38;2;154;148;143mL[38;2;129;115;96mv[38;2;150;124;98mX[38;2;153;117;73mv[38;2;120;88;56mj[38;2;78;60;52m_[38;2;164;149;129mL[38;2;240;227;206mM[38;2;193;180;156mw[38;2;176;163;134m0[38;2;251;236;191mM[38;2;252;236;186mM[38;2;254;237;202mW[38;2;255;239;212m&[38;2;255;240;215m&[38;2;254;242;220m8[38;2;254;244;219m8[38;2;255;246;218m8[38;2;247;239;209mW[38;2;230;213;174mh[38;2;250;225;181m*[38;2;251;225;172m*[38;2;252;224;168mo[38;2;252;224;172m*[38;2;253;227;174m*[38;2;252;226;173m*[38;2;252;225;174m*[38;2;252;226;179m*[38;2;254;233;192mM[38;2;244;227;188m*[38;2;219;199;159mb[38;2;223;199;155mb[38;2;236;209;150mk[38;2;205;169;98m0[38;2;196;146;70mU[38;2;178;124;64mz[38;2;81;44;24mi[38;2;37;22;19m,[38;2;59;48;33mi[38;2;100;81;55mt[38;2;109;85;56mf[38;2;81;62;40m_[38;2;26;20;12m\"[38;2;9;7;7m.[38;2;47;37;28ml[38;2;186;162;124m0[38;2;254;221;159mo[38;2;254;217;159ma[38;2;252;214;155ma[38;2;245;212;153mh[38;2;231;212;162mk[38;2;107;100;80mr[38;2;41;40;39ml[38;2;7;7;7m.[38;2;0;0;0m           [38;2;160;160;160mO[38;2;255;255;255m$$[38;2;247;254;254m@[38;2;210;140;143mO[38;2;253;0;8mj[38;2;255;1;12mj[38;2;255;2;12mj[38;2;255;1;11mj[38;2;255;0;4mf[38;2;210;111;114mC[38;2;242;250;250m@[38;2;255;255;255m$$[38;2;197;197;197mk[38;2;80;80;80mt[38;2;251;251;251m@[38;2;255;255;255m$$[38;2;239;240;239m8[38;2;225;81;88mY[38;2;255;0;3mf[38;2;255;0;11mj[38;2;255;0;10mj[38;2;255;0;9mj[38;2;248;0;7mf[38;2;194;113;117mJ[38;2;237;246;245m8[38;2;255;255;255m$$$[38;2;251;251;251m@@[38;2;252;253;252m$[38;2;255;255;255m$$$[38;2;217;221;219m*[38;2;203;55;63mu[38;2;249;0;2mf[38;2;249;0;7mf[38;2;248;0;8mf[38;2;249;0;8mf[38;2;240;0;8mt[38;2;217;145;149mm[38;2;249;253;254m$[38;2;249;255;254m$[38;2;199;148;151mZ[38;2;234;0;5mt[38;2;244;0;6mf[38;2;242;0;7mf[38;2;241;0;7mt[38;2;238;0;0mt[38;2;203;99;104mU[38;2;242;249;250m@[38;2;255;255;255m$$[38;2;233;241;241m8[38;2;200;72;78mc[38;2;236;0;0mt[38;2;235;0;7mt[38;2;234;0;6mt[38;2;233;0;6mt[38;2;234;0;6mt[38;2;233;0;3mt[38;2;231;0;0m1[38;2;229;0;0m1[38;2;228;0;0m1[38;2;227;0;0m1[38;2;226;0;0m11[38;2;224;0;1m11[38;2;222;0;0m1[38;2;224;0;0m1[38;2;200;15;23mt[38;2;213;206;207ma[38;2;255;255;255m$$$[38;2;64;64;64m-[38;2;0;0;0m");
  $display("[38;2;0;0;0m                           [38;2;5;5;3m [38;2;99;96;89mr[38;2;187;178;168mw[38;2;160;143;117mJ[38;2;131;106;79mn[38;2;119;89;57mj[38;2;131;101;77mn[38;2;228;207;174mh[38;2;255;248;215m8[38;2;189;178;159mw[38;2;119;106;89mn[38;2;246;233;193mM[38;2;249;236;188mM[38;2;254;238;203mW[38;2;255;239;214m&[38;2;255;240;215m&[38;2;255;241;219m8[38;2;255;244;219m8[38;2;255;246;219m8[38;2;251;240;211m&[38;2;235;217;184mo[38;2;251;229;189m#[38;2;252;228;183m#[38;2;252;229;183m#[38;2;253;232;189mM[38;2;254;236;195mM[38;2;254;236;199mW[38;2;255;237;203mW[38;2;255;238;209m&[38;2;254;240;212m&[38;2;254;241;214m&[38;2;253;242;218m&[38;2;253;243;221m8[38;2;255;247;221m8[38;2;255;244;213m&[38;2;253;229;183m#[38;2;254;207;137mk[38;2;241;179;103mw[38;2;177;129;79mY[38;2;86;63;39m_[38;2;38;27;18m,[38;2;35;23;20m,[38;2;20;10;7m'[38;2;46;32;24mI[38;2;123;98;76mx[38;2;208;178;125mm[38;2;247;217;149mh[38;2;251;221;161mo[38;2;253;225;173m*[38;2;252;222;168mo[38;2;252;220;170mo[38;2;212;191;145mq[38;2;149;140;102mY[38;2;45;43;33ml[38;2;0;0;0m            [38;2;158;158;158m0[38;2;255;255;255m$$[38;2;251;254;255m$[38;2;214;177;179md[38;2;205;68;73mc[38;2;202;61;67mv[38;2;203;62;68mv[38;2;202;61;67mv[38;2;206;62;68mv[38;2;211;156;159mw[38;2;248;251;251m@[38;2;255;255;255m$$[38;2;192;192;192mb[38;2;146;146;146mC[38;2;255;255;255m$$[38;2;254;255;255m$[38;2;224;202;204ma[38;2;205;71;78mc[38;2;201;58;65mu[38;2;200;59;67muu[38;2;202;58;65mu[38;2;199;91;97mY[38;2;218;217;216m*[38;2;253;255;255m$[38;2;255;255;255m$$[38;2;128;128;128mY[38;2;42;42;42m!![38;2;46;46;46mi[38;2;192;192;192mb[38;2;255;255;255m$$[38;2;249;253;252m@[38;2;203;178;179mp[38;2;200;68;73mv[38;2;196;58;64mu[38;2;195;58;65mu[38;2;194;58;65mn[38;2;196;57;62mn[38;2;199;104;109mU[38;2;237;237;239m&[38;2;252;255;255m$[38;2;208;182;184md[38;2;195;65;72mv[38;2;193;57;65mn[38;2;191;58;65mn[38;2;190;58;65mn[38;2;194;60;65mu[38;2;203;149;150mZ[38;2;248;250;251m@[38;2;255;255;255m$$[38;2;241;245;245mB[38;2;196;130;133mQ[38;2;190;58;63mn[38;2;187;58;64mn[38;2;186;58;64mn[38;2;186;58;63mnn[38;2;185;58;63mn[38;2;184;58;63mnn[38;2;184;57;63mn[38;2;183;58;63mn[38;2;182;58;64mnnnn[38;2;181;58;63mx[38;2;181;57;62mx[38;2;187;89;93mz[38;2;225;223;222m#[38;2;254;255;255m$[38;2;255;255;255m$$[38;2;62;62;62m_[38;2;0;0;0m");
  $display("[38;2;0;0;0m                           [38;2;21;21;12m^[38;2;139;133;78mc[38;2;141;124;83mc[38;2;200;183;152mw[38;2;162;146;114mJ[38;2;156;138;90mY[38;2;149;122;82mc[38;2;124;98;65mr[38;2;134;116;90mv[38;2;148;135;124mU[38;2;77;67;58m-[38;2;224;212;180mh[38;2;249;234;188m#[38;2;253;237;202mW[38;2;254;240;214m&[38;2;255;241;217m&[38;2;255;241;218m8[38;2;255;244;220m8[38;2;253;245;219m8[38;2;249;240;211mW[38;2;220;205;172mk[38;2;249;230;194mM[38;2;254;232;197mM[38;2;255;234;200mW[38;2;255;237;203mW[38;2;254;238;205mW[38;2;254;238;206mW[38;2;255;239;207mW[38;2;255;239;211m&[38;2;255;239;213m&[38;2;255;241;216m&[38;2;255;247;225m8[38;2;255;250;234mB[38;2;255;251;241m@[38;2;250;244;235mB[38;2;229;222;206m*[38;2;194;185;157mw[38;2;171;151;106mC[38;2;170;135;79mY[38;2;196;159;101mQ[38;2;178;144;99mJ[38;2;143;115;89mc[38;2;144;121;96mz[38;2;186;157;111mQ[38;2;248;214;152mh[38;2;249;214;144mh[38;2;250;217;148mh[38;2;252;223;165mo[38;2;251;224;172m*[38;2;251;224;170m*[38;2;249;221;171mo[38;2;193;175;136mZ[38;2;157;146;85mY[38;2;192;186;121mZ[38;2;52;52;34mi[38;2;0;0;0m           [38;2;65;65;65m-[38;2;236;236;236m&[38;2;255;255;255m$$[38;2;252;255;255m$[38;2;237;247;246mB[38;2;234;243;242m888[38;2;236;246;245m8[38;2;250;253;254m$[38;2;255;255;255m$$[38;2;249;249;249m@[38;2;92;92;92mr[38;2;53;53;53m~[38;2;233;233;233mW[38;2;255;255;255m$$[38;2;252;254;253m$[38;2;239;246;245mB[38;2;234;243;243m888[38;2;235;244;244m8[38;2;244;251;251m@[38;2;255;255;255m$$$[38;2;175;175;175mw[38;2;8;8;8m.[38;2;0;0;0m   [38;2;44;44;44m![38;2;223;223;223m#[38;2;255;255;255m$$$[38;2;239;248;248mB[38;2;235;243;243m8[38;2;234;243;243m8[38;2;234;243;242m8[38;2;235;244;243m8[38;2;243;248;248mB[38;2;255;255;255m$$[38;2;253;255;255m$[38;2;238;247;247mB[38;2;234;243;243m8[38;2;235;243;243m8[38;2;234;243;243m8[38;2;237;245;245m8[38;2;250;254;253m$[38;2;255;255;255m$$$$[38;2;247;253;252m@[38;2;236;244;244m8[38;2;234;243;243m8[38;2;235;243;243m88888888[38;2;235;243;244m8[38;2;235;243;243m8888[38;2;235;244;243m8[38;2;243;250;249m@[38;2;255;255;255m$$$[38;2;192;192;192mb[38;2;17;17;17m^[38;2;0;0;0m");
  $display("[38;2;0;0;0m                           [38;2;40;38;23mI[38;2;184;170;98mL[38;2;157;137;68mz[38;2;162;146;81mY[38;2;210;195;120mw[38;2;209;194;112mm[38;2;177;162;115mQ[38;2;168;157;132mQ[38;2;116;108;94mu[38;2;111;104;97mn[38;2;61;53;46m~[38;2;204;194;163mp[38;2;240;226;179m*[38;2;253;237;201mW[38;2;253;240;213m&[38;2;254;241;217m&[38;2;255;241;218m8[38;2;255;244;220m8[38;2;254;246;222m88[38;2;225;212;182ma[38;2;240;225;188m*[38;2;253;235;198mM[38;2;255;235;204mW[38;2;254;237;207mW[38;2;254;239;208mW[38;2;255;240;210m&[38;2;255;240;211m&[38;2;254;241;212m&[38;2;254;241;215m&[38;2;250;238;212mW[38;2;235;225;203m#[38;2;204;194;176md[38;2;169;157;137mQ[38;2;145;132;105mX[38;2;136;119;89mv[38;2;136;116;87mv[38;2;139;121;99mz[38;2;94;80;66mt[38;2;71;55;41m+[38;2;74;57;40m+[38;2;59;44;33m![38;2;63;49;44m~[38;2;85;68;48m-[38;2;147;126;94mz[38;2;234;213;162mh[38;2;250;228;169m*[38;2;250;225;170m*[38;2;252;225;170m*[38;2;250;223;170mo[38;2;251;228;188m#[38;2;167;151;129mL[38;2;79;68;41m_[38;2;178;172;97mL[38;2;134;132;85mc[38;2;0;0;0m            [38;2;42;42;42m![38;2;145;145;145mC[38;2;210;210;210ma[38;2;241;241;241m8[38;2;253;253;254m$[38;2;255;255;255m$$$[38;2;254;254;254m$[38;2;244;244;244mB[38;2;217;217;217m*[38;2;164;164;164mO[38;2;63;63;63m_[38;2;0;0;0m  [38;2;41;41;41ml[38;2;146;146;146mC[38;2;208;208;208ma[38;2;238;238;238m8[38;2;253;253;253m$[38;2;255;255;255m$$$$[38;2;250;250;250m@[38;2;231;231;231mW[38;2;188;188;188md[38;2;100;100;100mx[38;2;7;7;7m.[38;2;0;0;0m     [38;2;31;31;31m;[38;2;133;133;133mU[38;2;205;205;205mh[38;2;239;239;239m8[38;2;253;253;253m$[38;2;255;255;255m$$$[38;2;254;255;255m$[38;2;250;250;250m@[38;2;229;229;229mW[38;2;215;215;215m*[38;2;241;241;241m8[38;2;254;254;254m$[38;2;255;255;255m$$$[38;2;254;254;254m$[38;2;245;245;245mB[38;2;217;217;217m*[38;2;162;162;162mO[38;2;170;170;170mm[38;2;222;222;222m#[38;2;247;247;247m@[38;2;254;254;254m$[38;2;255;255;255m$$$$$$$$$$$$$$$[38;2;251;251;251m@[38;2;233;233;233mW[38;2;193;193;193mb[38;2;110;110;110mv[38;2;13;13;13m'[38;2;0;0;0m [38;2;0;0;0m");
  $display("[38;2;0;0;0m                          [38;2;7;8;5m.[38;2;89;86;58m1[38;2;168;157;97mJ[38;2;202;192;110mZ[38;2;221;206;101mw[38;2;201;178;84mQ[38;2;126;109;47mr[38;2;147;137;113mY[38;2;228;219;191mo[38;2;255;253;222mB[38;2;187;182;163mw[38;2;35;29;22m;[38;2;179;171;148mZ[38;2;240;230;186m*[38;2;251;238;199mW[38;2;253;238;211m&[38;2;255;240;216m&[38;2;255;241;218m8[38;2;254;243;219m8[38;2;254;244;219m8[38;2;255;244;226m8[38;2;236;224;201m#[38;2;228;215;181ma[38;2;252;237;200mW[38;2;254;236;204mW[38;2;255;238;208mW[38;2;255;240;209m&[38;2;255;241;210m&[38;2;254;239;211m&[38;2;250;238;209mW[38;2;201;188;162mp[38;2;150;135;110mY[38;2;125;110;82mn[38;2;130;116;87mv[38;2;169;154;124mL[38;2;201;186;157mq[38;2;222;209;182mh[38;2;240;229;205mM[38;2;253;245;223m8[38;2;243;233;214mW[38;2;203;193;175md[38;2;160;152;136mL[38;2;155;148;129mC[38;2;211;201;183mk[38;2;190;178;160mw[38;2;115;99;82mx[38;2;136;119;90mc[38;2;231;211;170mh[38;2;251;231;182m#[38;2;251;228;177m*[38;2;252;227;181m#[38;2;228;210;175mh[38;2;117;101;71mx[38;2;122;114;68mn[38;2;164;163;100mC[38;2;75;75;52m-[38;2;0;0;0m              [38;2;5;5;5m.[38;2;30;30;30m;[38;2;47;47;47mi[38;2;49;49;49mi[38;2;48;48;48mi[38;2;49;49;49mi[38;2;48;48;48mi[38;2;34;34;34mI[38;2;9;9;9m.[38;2;0;0;0m      [38;2;4;4;4m [38;2;27;27;27m,[38;2;46;46;46mi[38;2;49;49;49mi[38;2;48;48;48mii[38;2;49;49;49mi[38;2;42;42;42m![38;2;19;19;19m\"[38;2;0;0;0m          [38;2;3;3;3m [38;2;27;27;27m,[38;2;46;46;46mi[38;2;49;49;49mi[38;2;48;48;48mii[38;2;49;49;49mi[38;2;43;43;43m![38;2;19;19;19m\"[38;2;7;7;7m.[38;2;30;30;30m;[38;2;47;47;47mi[38;2;49;49;49mi[38;2;48;48;48mi[38;2;49;49;49mi[38;2;48;48;48mi[38;2;35;35;35mI[38;2;9;9;9m.[38;2;0;0;0m  [38;2;13;13;13m'[38;2;38;38;38ml[38;2;48;48;48mi[38;2;49;49;49mi[38;2;48;48;48miiiiiiiiiiiii[38;2;49;49;49mi[38;2;44;44;44m![38;2;21;21;21m\"[38;2;0;0;0m    [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;5;5;3m [38;2;119;120;85mu[38;2;194;189;118mZ[38;2;197;186;107mO[38;2;171;162;83mJ[38;2;222;198;101mm[38;2;166;133;56mc[38;2;122;96;46mj[38;2;149;131;78mz[38;2;153;136;83mX[38;2;136;121;94mc[38;2;81;75;65m?[38;2;8;5;4m.[38;2;139;130;113mX[38;2;242;231;194m#[38;2;250;236;198mM[38;2;251;236;207mW[38;2;255;239;216m&[38;2;255;242;218m8[38;2;254;242;218m8[38;2;253;241;216m&[38;2;254;241;222m8[38;2;250;238;218m&[38;2;227;216;185ma[38;2;249;236;201mM[38;2;254;237;210mW[38;2;255;238;212m&[38;2;255;240;213m&[38;2;255;241;213m&[38;2;254;242;213m&[38;2;250;238;208mW[38;2;200;184;151mw[38;2;189;173;135mZ[38;2;229;213;175mh[38;2;252;236;202mW[38;2;247;233;201mM[38;2;249;236;208mW[38;2;255;249;223m8[38;2;255;248;224m8[38;2;255;248;221m8[38;2;255;246;214m8[38;2;255;246;211m&[38;2;255;247;210m&[38;2;255;245;207m&[38;2;255;239;198mW[38;2;255;244;198mW[38;2;235;214;171ma[38;2;158;133;100mY[38;2;206;181;144mw[38;2;253;230;182m#[38;2;251;228;178m*[38;2;252;235;189mM[38;2;147;138;110mY[38;2;105;89;54mt[38;2;131;122;74mu[38;2;47;47;31ml[38;2;0;0;0m                                                                                             [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;31;30;24m;[38;2;187;186;135mZ[38;2;191;183;89mQ[38;2;223;210;95mw[38;2;202;194;97mO[38;2;166;153;73mY[38;2;206;188;87mO[38;2;196;176;75mL[38;2;185;165;82mC[38;2;207;187;133mw[38;2;198;184;154mw[38;2;59;52;46m~[38;2;0;0;0m [38;2;75;66;58m-[38;2;240;226;197m#[38;2;251;236;200mW[38;2;252;237;204mW[38;2;254;240;215m&[38;2;254;242;218m8[38;2;254;243;218m8[38;2;254;242;217m&[38;2;254;242;218m8[38;2;255;243;222m8[38;2;247;235;208mW[38;2;248;233;204mM[38;2;253;237;211mW[38;2;255;238;212m&[38;2;255;240;214m&[38;2;255;241;214m&[38;2;254;243;215m&[38;2;253;243;212m&[38;2;247;227;184m*[38;2;240;217;169ma[38;2;180;159;127mQ[38;2;190;173;144mZ[38;2;226;210;175mh[38;2;232;215;176ma[38;2;227;209;170mh[38;2;224;205;167mk[38;2;226;202;162mb[38;2;227;202;157mb[38;2;226;199;151mb[38;2;227;197;147md[38;2;228;196;143md[38;2;217;186;136mq[38;2;191;163;115m0[38;2;177;150;100mC[38;2;231;202;146mb[38;2;250;221;163mo[38;2;251;221;166mo[38;2;253;225;174m*[38;2;234;222;184mo[38;2;65;59;48m+[38;2;84;71;49m-[38;2;106;96;74mr[38;2;16;14;14m^[38;2;0;0;0m                                                                                             [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;27;26;20m,[38;2;125;119;69mn[38;2;206;190;90mO[38;2;193;172;61mC[38;2;250;239;135ma[38;2;228;217;115mp[38;2;204;187;83m0[38;2;157;143;71mz[38;2;168;156;123mL[38;2;251;236;207mW[38;2;255;246;213m8[38;2;150;141;128mJ[38;2;0;0;0m [38;2;46;41;38ml[38;2;238;224;198m#[38;2;253;237;199mW[38;2;253;237;203mW[38;2;254;240;215m&[38;2;253;241;220m8[38;2;255;243;221m88[38;2;255;243;220m8[38;2;255;244;221m8[38;2;239;226;203m#[38;2;230;215;192mo[38;2;253;239;214m&[38;2;253;240;214m&[38;2;255;242;216m&[38;2;254;242;218m8[38;2;253;244;223m8[38;2;254;244;225m8[38;2;251;235;203mW[38;2;230;206;165mk[38;2;103;80;60mt[38;2;30;15;11m^[38;2;29;20;16m\"[38;2;37;30;22m;[38;2;37;28;21m;[38;2;43;35;27mI[38;2;44;36;28mI[38;2;45;34;26mI[38;2;43;31;24mI[38;2;42;29;20m;[38;2;39;26;18m,[38;2;32;19;13m\"[38;2;43;27;19m;[38;2;107;86;62mf[38;2;220;194;147mp[38;2;250;222;162mo[38;2;250;219;165mo[38;2;255;227;182m#[38;2;192;180;154mw[38;2;54;51;41mi[38;2;93;83;58mt[38;2;104;98;74mr[38;2;7;7;6m.[38;2;0;0;0m                   [38;2;0;0;1m [38;2;0;0;0m    [38;2;0;0;1m [38;2;0;0;0m [38;2;5;5;7m.[38;2;10;10;10m'[38;2;14;14;13m'[38;2;40;40;38ml[38;2;83;83;79mt[38;2;108;108;102mu[38;2;93;93;88mj[38;2;39;38;37ml[38;2;5;5;5m.[38;2;0;0;0m                                                          [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;16;16;9m'[38;2;164;157;81mU[38;2;210;189;79m0[38;2;179;162;57mY[38;2;251;241;137ma[38;2;224;208;108mq[38;2;229;204;90mw[38;2;164;148;77mY[38;2;166;159;137mQ[38;2;237;224;197m*[38;2;255;241;213m&[38;2;198;190;173mp[38;2;9;8;7m.[38;2;30;27;23m,[38;2;207;199;173mb[38;2;252;239;203mW[38;2;252;237;203mW[38;2;254;239;212m&[38;2;255;241;217m&[38;2;255;244;220m8[38;2;255;244;222m8[38;2;255;242;223m8[38;2;255;243;225m8[38;2;241;230;211mM[38;2;229;219;199m*[38;2;254;244;224m8[38;2;253;243;223m8[38;2;254;244;224m8[38;2;253;245;225m8[38;2;253;246;226m8[38;2;255;246;227m8[38;2;255;246;226m8[38;2;254;241;215m&[38;2;237;224;191m*[38;2;197;187;159mq[38;2;155;148;125mC[38;2;157;150;125mC[38;2;187;175;146mZ[38;2;206;188;154mq[38;2;212;190;151mp[38;2;211;185;148mq[38;2;203;173;137mm[38;2;182;146;105mC[38;2;179;141;92mU[38;2;183;148;100mC[38;2;185;156;106mL[38;2;235;203;154mk[38;2;254;221;168mo[38;2;251;219;162ma[38;2;248;220;172mo[38;2;247;225;195m#[38;2;110;102;89mx[38;2;47;48;36m![38;2;74;68;44m_[38;2;78;76;56m?[38;2;0;0;0m                    [38;2;1;0;1m [38;2;75;72;64m?[38;2;165;160;136mQ[38;2;143;136;116mY[38;2;109;101;90mx[38;2;140;133;125mY[38;2;178;171;164mm[38;2;200;195;182mb[38;2;210;205;187mk[38;2;205;197;178mb[38;2;170;162;140m0[38;2;233;226;202m#[38;2;255;255;231m@[38;2;235;229;208mM[38;2;145;141;125mU[38;2;87;83;70mt[38;2;119;116;107mv[38;2;66;65;58m_[38;2;17;17;16m^[38;2;0;0;0m                                                       [38;2;0;0;0m");
  $display("[38;2;0;0;0m                         [38;2;24;24;16m\"[38;2;196;188;121mZ[38;2;194;176;75mL[38;2;187;172;65mJ[38;2;245;235;131mh[38;2;198;180;93m0[38;2;205;180;77mQ[38;2;162;147;81mY[38;2;191;187;166mq[38;2;235;226;198m*[38;2;253;240;214m&[38;2;244;236;216mW[38;2;75;71;65m?[38;2;0;0;0m [38;2;142;140;117mU[38;2;239;231;196m#[38;2;255;244;207m&[38;2;254;241;204mW[38;2;254;239;206mW[38;2;255;241;211m&[38;2;255;243;220m8[38;2;254;244;226m8[38;2;254;246;228m8[38;2;242;235;217mW[38;2;232;225;207m#[38;2;255;249;230mB[38;2;254;247;228mB[38;2;254;246;228m88[38;2;254;246;227m8[38;2;255;246;227m8[38;2;255;246;230mB[38;2;255;246;229mB[38;2;255;249;227mB[38;2;255;251;227mB[38;2;255;253;228mB[38;2;255;252;224mB[38;2;255;243;210m&[38;2;248;229;187m#[38;2;251;228;177m*[38;2;255;231;185m#[38;2;200;164;123mO[38;2;209;166;109mO[38;2;250;204;128mb[38;2;253;205;134mk[38;2;250;211;144mk[38;2;252;217;150ma[38;2;253;217;152ma[38;2;249;218;157ma[38;2;250;230;188m#[38;2;189;176;154mm[38;2;95;84;71mf[38;2;64;58;50m+[38;2;65;63;47m+[38;2;51;52;42mi[38;2;0;0;0m                    [38;2;20;17;16m^[38;2;202;189;166mp[38;2;255;243;193mW[38;2;255;237;187mM[38;2;252;230;186m#[38;2;224;208;171mk[38;2;214;203;174mk[38;2;241;231;203mM[38;2;252;241;207mW[38;2;243;227;194m#[38;2;213;195;162md[38;2;164;146;113mJ[38;2;206;190;158mp[38;2;215;203;169mb[38;2;234;222;188mo[38;2;157;140;111mU[38;2;197;183;154mw[38;2;251;242;208mW[38;2;219;212;184mh[38;2;135;133;118mY[38;2;41;42;38ml[38;2;17;17;17m^[38;2;0;0;0m       [38;2;1;1;2m [38;2;5;4;5m [38;2;0;0;0m                                           [38;2;0;0;0m");
  $display("[38;2;0;0;0m                    [38;2;1;2;3m [38;2;6;6;7m.[38;2;0;0;0m   [38;2;17;17;15m^[38;2;173;169;113mQ[38;2;186;170;73mC[38;2;187;171;65mJ[38;2;243;234;132mh[38;2;172;154;78mU[38;2;175;152;60mY[38;2;151;139;80mz[38;2;193;189;168mp[38;2;238;228;200m#[38;2;253;238;214m&[38;2;255;245;222m8[38;2;218;212;192ma[38;2;97;94;82mj[38;2;49;43;37m![38;2;92;85;74mf[38;2;175;167;147mO[38;2;231;223;189mo[38;2;252;240;197mW[38;2;255;238;196mW[38;2;252;237;204mW[38;2;252;241;213m&[38;2;247;241;218m&[38;2;237;231;208mM[38;2;220;211;189ma[38;2;237;227;206m#[38;2;248;238;217m&[38;2;254;245;227m8[38;2;254;245;228m8[38;2;254;245;227m8[38;2;254;246;226m8[38;2;253;245;225m8[38;2;253;245;223m8[38;2;253;246;220m8[38;2;254;246;221m8[38;2;255;243;221m8[38;2;255;242;211m&[38;2;250;233;194mM[38;2;243;225;179m*[38;2;248;228;178m*[38;2;240;217;173ma[38;2;175;147;115mC[38;2;136;106;67mn[38;2;204;171;108mO[38;2;245;208;138mk[38;2;247;212;149mh[38;2;252;218;157ma[38;2;252;219;156ma[38;2;250;225;176m*[38;2;244;231;205mM[38;2;139;130;108mX[38;2;157;145;114mJ[38;2;78;65;47m_[38;2;49;49;42mi[38;2;18;20;18m^[38;2;0;0;0m                    [38;2;13;13;11m'[38;2;161;149;130mC[38;2;252;229;184m#[38;2;255;233;174m#[38;2;255;232;174m#[38;2;254;228;172m*[38;2;247;222;174mo[38;2;220;194;150md[38;2;180;152;106mC[38;2;169;138;91mY[38;2;160;129;84mX[38;2;138;107;68mn[38;2;111;88;50mf[38;2;117;95;54mj[38;2;159;134;93mY[38;2;171;147;112mC[38;2;128;114;85mu[38;2;203;192;168mp[38;2;210;198;174mb[38;2;182;172;154mZ[38;2;108;103;92mn[38;2;95;94;87mr[38;2;74;73;68m?[38;2;71;68;64m-[38;2;82;80;72mt[38;2;95;92;83mj[38;2;89;86;77mf[38;2;123;119;110mc[38;2;156;151;139mL[38;2;184;179;162mw[38;2;196;191;177md[38;2;89;86;80mf[38;2;6;6;5m.[38;2;0;0;0m                                         [38;2;0;0;0m");
  $display("[38;2;0;0;0m               [38;2;0;0;2m [38;2;40;41;37ml[38;2;94;92;69mf[38;2;132;128;84mv[38;2;158;154;93mU[38;2;186;182;106m0[38;2;197;191;105mO[38;2;159;155;83mY[38;2;49;50;29m![38;2;1;1;3m [38;2;9;10;9m.[38;2;162;159;105mC[38;2;188;174;81mL[38;2;173;156;57mY[38;2;232;222;128mb[38;2;149;134;59mv[38;2;155;138;49mv[38;2;120;109;56mr[38;2;186;179;159mw[38;2;239;224;197m#[38;2;254;239;212m&[38;2;252;238;216m&[38;2;255;245;219m8[38;2;253;246;217m8[38;2;205;198;176mb[38;2;110;105;92mn[38;2;35;29;26m;[38;2;40;34;30mI[38;2;125;117;104mc[38;2;192;177;151mm[38;2;204;190;152mq[38;2;206;193;151mp[38;2;209;195;162md[38;2;204;189;162mp[38;2;208;193;165md[38;2;245;231;204mM[38;2;253;241;217m&[38;2;253;244;219m8[38;2;255;245;221m8[38;2;255;245;224m8[38;2;254;244;222m8[38;2;254;244;219m8[38;2;254;245;218m8[38;2;253;245;217m8[38;2;255;243;218m8[38;2;255;240;212m&[38;2;251;234;199mM[38;2;249;229;185m#[38;2;250;228;184m#[38;2;198;179;137mm[38;2;150;131;101mX[38;2;95;81;65mt[38;2;40;25;13m,[38;2;191;167;125mO[38;2;254;223;157mo[38;2;253;222;157ma[38;2;253;220;158ma[38;2;248;221;164mo[38;2;255;241;204mW[38;2;175;165;153mO[38;2;130;121;96mc[38;2;241;223;180mo[38;2;133;119;94mc[38;2;18;16;14m^[38;2;3;3;4m [38;2;0;0;0m                     [38;2;16;13;11m'[38;2;109;97;84mx[38;2;177;162;128mQ[38;2;215;194;150mp[38;2;216;189;138mq[38;2;221;190;129mq[38;2;228;195;128mp[38;2;220;185;114mm[38;2;218;182;110mm[38;2;209;172;108mO[38;2;193;153;106mL[38;2;155;127;94mX[38;2;130;111;88mu[38;2;129;114;95mv[38;2;160;149;131mC[38;2;196;188;169mp[38;2;220;210;190ma[38;2;234;221;201m*[38;2;235;223;202m#[38;2;186;175;153mm[38;2;131;124;106mz[38;2;113;106;98mn[38;2;224;216;201mo[38;2;255;249;215m8[38;2;255;249;216m8[38;2;233;222;192m*[38;2;169;157;130mQ[38;2;255;244;211m&[38;2;255;247;206m&[38;2;255;250;208m&[38;2;229;224;195m*[38;2;63;62;53m+[38;2;0;0;0m                                         [38;2;0;0;0m");
  $display("[38;2;0;0;0m           [38;2;0;0;1m [38;2;0;0;0m  [38;2;53;53;48m~[38;2;71;67;48m_[38;2;204;198;148mp[38;2;255;253;172mM[38;2;255;246;143mo[38;2;255;242;117mh[38;2;255;240;104mk[38;2;254;237;95mb[38;2;240;224;93mp[38;2;205;193;101mZ[38;2;60;56;38m~[38;2;47;49;46mi[38;2;161;159;106mC[38;2;158;140;71mz[38;2;155;131;58mv[38;2;195;179;101m0[38;2;136;121;56mn[38;2;149;132;56mv[38;2;95;86;46m1[38;2;191;185;165mq[38;2;236;221;195m*[38;2;254;239;210m&[38;2;252;239;211m&[38;2;252;240;212m&[38;2;253;241;212m&[38;2;255;242;213m&[38;2;255;245;213m&[38;2;216;206;178mk[38;2;105;99;84mx[38;2;16;13;8m'[38;2;16;10;10m'[38;2;46;40;33ml[38;2;95;87;70mf[38;2;137;125;97mz[38;2;202;189;151mq[38;2;215;201;160mb[38;2;215;201;166mb[38;2;239;227;196m#[38;2;250;243;207mW[38;2;252;244;215m&[38;2;254;244;218m8[38;2;254;243;216m&[38;2;255;243;214m&[38;2;254;241;211m&[38;2;253;238;208mW[38;2;255;238;210m&[38;2;254;237;204mW[38;2;240;224;188m*[38;2;209;194;164md[38;2;145;131;112mY[38;2;57;46;39mi[38;2;43;34;31mI[38;2;31;24;23m,[38;2;32;20;19m,[38;2;100;85;66mf[38;2;173;150;109mC[38;2;238;204;150mk[38;2;250;222;164mo[38;2;248;236;197mM[38;2;239;239;222mW[38;2;62;55;52m+[38;2;156;140;111mU[38;2;222;200;155mb[38;2;135;123;100mz[38;2;19;17;17m^[38;2;0;0;1m [38;2;0;0;0m                        [38;2;12;10;9m'[38;2;27;21;17m\"[38;2;49;42;29ml[38;2;61;53;36mi[38;2;60;51;35mi[38;2;65;55;39m~[38;2;121;108;88mn[38;2;147;129;107mX[38;2;145;129;107mX[38;2;196;182;158mw[38;2;242;228;196m#[38;2;255;237;200mW[38;2;255;240;197mW[38;2;255;239;192mM[38;2;254;238;188mM[38;2;254;237;189mM[38;2;255;242;198mW[38;2;236;221;182mo[38;2;152;136;115mU[38;2;148;134;114mY[38;2;241;228;191m#[38;2;231;217;177ma[38;2;242;226;192m#[38;2;187;169;140mZ[38;2;190;173;135mZ[38;2;216;200;156md[38;2;205;193;148mq[38;2;200;189;157mq[38;2;80;78;67m1[38;2;0;0;0m    [38;2;0;0;1m [38;2;5;4;5m [38;2;5;6;6m.[38;2;10;10;11m'[38;2;0;0;0m                                 [38;2;0;0;0m");
  $display("[38;2;0;0;0m            [38;2;11;11;9m'[38;2;117;111;78mn[38;2;231;215;135mb[38;2;224;204;102mw[38;2;209;193;92mO[38;2;218;204;108mw[38;2;250;234;123mh[38;2;251;232;99mb[38;2;252;229;89md[38;2;253;232;93mb[38;2;197;177;76mL[38;2;207;182;92mO[38;2;143;131;80mc[38;2;51;53;46mi[38;2;148;148;96mY[38;2;144;127;64mv[38;2;142;118;57mn[38;2;167;149;83mU[38;2;136;120;62mu[38;2;146;130;64mv[38;2;77;69;39m_[38;2;187;182;166mw[38;2;240;228;199m#[38;2;255;240;211m&[38;2;255;239;210m&[38;2;255;241;211m&[38;2;255;239;211m&[38;2;255;235;207mW[38;2;255;233;196mM[38;2;255;237;193mM[38;2;249;232;189m#[38;2;195;182;148mw[38;2;96;87;73mf[38;2;21;18;15m^[38;2;0;0;0m [38;2;18;14;13m^[38;2;82;76;62m?[38;2;146;138;109mY[38;2;188;176;142mZ[38;2;214;200;166mb[38;2;253;241;206mW[38;2;255;244;215m8[38;2;255;241;213m&[38;2;255;239;209m&[38;2;255;238;204mW[38;2;255;240;203mW[38;2;253;236;203mW[38;2;207;190;168md[38;2;139;126;111mX[38;2;77;69;60m-[38;2;40;33;27mI[38;2;35;28;23m;[38;2;41;31;25mI[38;2;51;35;25ml[38;2;55;36;22ml[38;2;65;46;31mi[38;2;45;29;19m;[38;2;29;13;9m^[38;2;98;79;62mt[38;2;193;179;148mm[38;2;255;255;238m@[38;2;174;172;167mm[38;2;52;45;37m![38;2;186;174;138mZ[38;2;183;166;127m0[38;2;126;117;97mv[38;2;12;12;13m'[38;2;0;0;0m                       [38;2;17;17;12m^[38;2;41;41;30ml[38;2;58;58;46m~[38;2;26;25;20m,[38;2;6;5;5m.[38;2;33;33;35mI[38;2;94;93;93mr[38;2;163;162;154m0[38;2;235;231;216mM[38;2;238;232;211mM[38;2;157;147;130mC[38;2;145;130;105mX[38;2;176;159;116mL[38;2;236;215;165mh[38;2;234;213;163mh[38;2;226;204;154mb[38;2;223;200;149md[38;2;222;197;150md[38;2;217;192;150mp[38;2;211;187;147mq[38;2;201;180;142mw[38;2;181;166;132m0[38;2;182;170;141mO[38;2;135;124;102mz[38;2;140;127;110mX[38;2;172;154;131mQ[38;2;200;179;144mw[38;2;178;160;119mQ[38;2;172;155;117mL[38;2;194;179;145mm[38;2;185;174;150mZ[38;2;171;162;145m0[38;2;171;159;146m0[38;2;169;160;144m0[38;2;163;157;143mQ[38;2;120;114;104mv[38;2;153;149;141mL[38;2;196;194;183md[38;2;206;205;192mk[38;2;163;163;155mO[38;2;50;51;48mi[38;2;0;0;0m                               [38;2;0;0;0m");
  $display("[38;2;0;0;0m          [38;2;3;3;4m [38;2;63;64;43m+[38;2;179;174;107mQ[38;2;247;226;122mk[38;2;247;218;90mp[38;2;247;218;87mp[38;2;247;217;95mp[38;2;208;182;73mQ[38;2;232;210;100mq[38;2;254;233;100mb[38;2;252;231;88md[38;2;246;229;98md[38;2;139;122;57mu[38;2;198;173;95mQ[38;2;169;151;85mU[38;2;0;0;0m [38;2;137;134;86mz[38;2;167;151;80mY[38;2;144;121;63mu[38;2;148;126;75mc[38;2;137;118;64mu[38;2;108;94;45mt[38;2;56;45;23ml[38;2;176;170;155mZ[38;2;229;218;188mo[38;2;253;238;208mW[38;2;254;238;209mW[38;2;254;240;210m&[38;2;254;238;208mW[38;2;254;235;203mW[38;2;254;233;193mM[38;2;254;232;184m#[38;2;251;229;178m*[38;2;247;226;177m*[38;2;206;189;147mq[38;2;119;107;82mn[38;2;27;20;14m\"[38;2;8;6;8m.[38;2;0;0;0m [38;2;7;6;4m.[38;2;51;48;41mi[38;2;120;113;94mu[38;2;201;190;165mp[38;2;229;215;184ma[38;2;237;222;185mo[38;2;231;217;179ma[38;2;213;200;167mb[38;2;189;179;152mm[38;2;108;98;83mx[38;2;60;51;42m~[38;2;66;56;45m+[38;2;79;67;54m-[38;2;81;66;51m-[38;2;96;79;60mt[38;2;101;76;55m1[38;2;101;69;43m?[38;2;111;74;44m1[38;2;118;76;46mt[38;2;138;91;62mx[38;2;110;77;50mt[38;2;62;45;32mi[38;2;54;48;40mi[38;2;148;147;139mC[38;2;70;65;60m-[38;2;84;73;58m?[38;2;166;155;126mL[38;2;237;226;200m#[38;2;173;167;154mO[38;2;10;11;12m'[38;2;0;0;0m                   [38;2;0;1;2m [38;2;38;38;32mI[38;2;101;101;76mr[38;2;154;153;106mU[38;2;180;176;127mO[38;2;186;182;130mZ[38;2;188;186;139mm[38;2;173;170;142mO[38;2;184;179;165mw[38;2;196;189;178mp[38;2;178;169;154mZ[38;2;186;176;151mm[38;2;197;190;168mp[38;2;172;164;148mO[38;2;144;131;117mY[38;2;149;133;107mY[38;2;184;166;126m0[38;2;193;171;127mOO[38;2;198;172;131mZ[38;2;205;175;136mm[38;2;210;178;139mw[38;2;216;187;145mq[38;2;230;206;161mk[38;2;237;216;174ma[38;2;223;204;169mk[38;2;194;179;151mw[38;2;137;123;99mz[38;2;160;145;119mJ[38;2;238;218;174ma[38;2;253;229;178m#[38;2;235;218;173ma[38;2;188;176;137mZ[38;2;168;158;125mL[38;2;224;211;181mh[38;2;255;246;216m8[38;2;255;244;214m&&[38;2;255;247;221m8[38;2;231;223;201m*[38;2;154;148;130mC[38;2;229;224;205m*[38;2;255;254;233m@[38;2;255;255;242m@[38;2;187;189;183mp[38;2;8;9;10m.[38;2;0;0;0m                              [38;2;0;0;0m");
  $display("[38;2;0;0;0m       [38;2;7;8;10m.[38;2;31;32;26m;[38;2;73;69;46m_[38;2;170;158;100mC[38;2;236;220;117md[38;2;246;224;97md[38;2;243;214;86mq[38;2;244;215;86mq[38;2;245;216;83mq[38;2;249;218;86mp[38;2;222;193;80mZ[38;2;218;193;81mO[38;2;254;235;96mb[38;2;250;232;99mb[38;2;160;149;74mX[38;2;69;54;25mi[38;2;231;208;114mp[38;2;150;132;66mc[38;2;22;19;10m^[38;2;134;127;92mc[38;2;189;175;95mQ[38;2;154;135;63mc[38;2;139;116;67mu[38;2;128;108;61mx[38;2;109;94;52mf[38;2;49;40;21mI[38;2;173;169;160mZ[38;2;212;204;180mk[38;2;249;234;202mM[38;2;253;238;209mW[38;2;254;238;207mW[38;2;254;238;203mW[38;2;254;236;201mW[38;2;253;234;192mM[38;2;254;232;184m#[38;2;250;226;172m*[38;2;244;218;160ma[38;2;247;219;163ma[38;2;231;210;166mh[38;2;159;145;118mJ[38;2;68;61;51m_[38;2;16;12;10m'[38;2;1;0;0m [38;2;0;0;0m  [38;2;26;23;19m\"[38;2;74;67;58m-[38;2;121;110;97mu[38;2;103;94;77mj[38;2;77;69;59m-[38;2;40;30;24m;[38;2;78;65;51m-[38;2;114;102;77mx[38;2;109;92;67mj[38;2;100;79;54m1[38;2;95;74;53m1[38;2;84;62;44m_[38;2;85;61;46m-[38;2;67;45;34mi[38;2;59;38;32m![38;2;56;33;28ml[38;2;65;40;27m![38;2;65;43;28m![38;2;83;67;49m-[38;2;44;40;31ml[38;2;0;0;0m [38;2;33;30;22m;[38;2;144;130;111mY[38;2;162;148;130mC[38;2;254;248;235mB[38;2;175;170;163mZ[38;2;9;11;11m'[38;2;0;0;0m                [38;2;10;11;10m'[38;2;32;33;25m;[38;2;95;94;64mf[38;2;171;172;113mQ[38;2;193;192;131mm[38;2;185;183;141mZ[38;2;195;193;165mp[38;2;188;185;171mq[38;2;180;176;165mm[38;2;180;175;163mm[38;2;164;157;150m0[38;2;130;121;113mz[38;2;127;117;96mv[38;2;187;173;140mZ[38;2;225;210;175mh[38;2;185;175;151mm[38;2;119;112;97mu[38;2;144;136;119mU[38;2;145;137;110mY[38;2;189;176;141mZ[38;2;246;229;186m#[38;2;250;227;181m*[38;2;252;226;182m#[38;2;255;226;181m#[38;2;253;224;179m*[38;2;238;213;169ma[38;2;202;180;143mw[38;2;180;158;127mQ[38;2;171;146;116mC[38;2;201;177;137mm[38;2;236;209;164mh[38;2;251;223;173m*[38;2;246;221;166mo[38;2;248;229;186m#[38;2;247;240;210mW[38;2;237;234;213mM[38;2;161;153;135mL[38;2;164;152;131mL[38;2;203;188;162mp[38;2;220;203;172mk[38;2;228;211;179ma[38;2;222;205;176mk[38;2;208;196;168md[38;2;162;154;127mL[38;2;181;177;150mZ[38;2;232;230;210mM[38;2;205;205;194mk[38;2;74;75;76m1[38;2;1;1;2m [38;2;0;0;0m                              [38;2;0;0;0m");
  $display("[38;2;0;0;0m    [38;2;0;0;1m [38;2;28;31;26m;[38;2;80;82;64m1[38;2;136;133;89mz[38;2;198;186;111mZ[38;2;247;224;117mb[38;2;255;223;100mb[38;2;246;213;86mq[38;2;244;214;86mq[38;2;244;215;85mq[38;2;245;216;85mq[38;2;247;217;85mp[38;2;243;215;90mq[38;2;212;189;82mO[38;2;235;213;97mq[38;2;253;233;90mb[38;2;228;210;102mq[38;2;56;47;24m![38;2;129;114;64mn[38;2;243;221;113mb[38;2;117;105;53mj[38;2;25;23;14m\"[38;2;89;83;58m1[38;2;186;174;101mQ[38;2;152;134;58mv[38;2;140;116;60mn[38;2;112;89;44mt[38;2;130;113;62mn[38;2;65;57;29mi[38;2;174;172;165mm[38;2;225;218;200mo[38;2;244;228;199m#[38;2;255;238;206mW[38;2;255;240;206mW[38;2;255;240;202mW[38;2;255;238;195mW[38;2;252;233;185m#[38;2;253;229;178m#[38;2;252;224;171m*[38;2;247;217;163ma[38;2;243;217;161ma[38;2;246;229;190m#[38;2;255;247;222m8[38;2;175;168;152mZ[38;2;74;69;56m-[38;2;31;26;19m,[38;2;3;0;0m [38;2;0;0;0m   [38;2;2;0;0m [38;2;3;0;0m [38;2;26;21;18m\"[38;2;88;78;66m1[38;2;111;96;72mr[38;2;98;83;54mt[38;2;103;83;58mt[38;2;99;77;53m1[38;2;93;70;48m?[38;2;96;73;54m1[38;2;81;62;47m_[38;2;54;40;30ml[38;2;55;45;37m![38;2;65;56;49m+[38;2;37;30;24m;[38;2;24;20;17m\"[38;2;8;6;5m.[38;2;0;0;0m  [38;2;47;44;35m![38;2;204;188;163mp[38;2;180;160;138m0[38;2;216;200;179mk[38;2;126;117;106mc[38;2;6;7;8m.[38;2;7;8;7m.[38;2;2;3;4m [38;2;0;0;1m [38;2;0;0;0m        [38;2;14;12;11m'[38;2;37;35;23m;[38;2;75;73;42m_[38;2;127;124;77mu[38;2;177;169;108mQ[38;2;206;197;118mm[38;2;224;218;113mp[38;2;232;222;118md[38;2;198;186;117mZ[38;2;160;151;121mC[38;2;206;202;193mk[38;2;212;212;209mo[38;2;197;194;182md[38;2;188;183;170mq[38;2;177;168;153mZ[38;2;185;173;149mZ[38;2;211;195;160md[38;2;232;216;174ma[38;2;206;189;151mq[38;2;167;152;120mC[38;2;205;194;175md[38;2;252;244;228m8[38;2;241;234;216mW[38;2;201;196;176md[38;2;126;117;102mc[38;2;177;166;147mO[38;2;242;230;203mM[38;2;230;218;190mo[38;2;192;179;151mw[38;2;165;150;127mL[38;2;111;95;79mr[38;2;113;95;80mx[38;2;189;169;136mO[38;2;236;215;166mh[38;2;247;226;176m*[38;2;249;229;185m#[38;2;253;236;200mW[38;2;250;240;210mW[38;2;233;228;202m#[38;2;219;210;178mh[38;2;217;200;157md[38;2;217;195;154md[38;2;189;167;137mO[38;2;153;130;96mX[38;2;234;214;168mh[38;2;233;213;166mh[38;2;231;210;165mh[38;2;222;202;157mb[38;2;216;198;160md[38;2;186;172;145mZ[38;2;119;113;98mv[38;2;43;43;40m![38;2;0;0;0m [38;2;0;0;1m [38;2;0;0;0m                              [38;2;0;0;0m");
  $display("[38;2;0;0;0m  [38;2;25;25;20m,[38;2;79;77;50m-[38;2;132;127;80mv[38;2;193;185;115mO[38;2;225;214;116mp[38;2;244;224;104md[38;2;251;222;91md[38;2;249;216;85mp[38;2;249;214;88mp[38;2;248;215;87mp[38;2;246;216;86mq[38;2;247;216;85mq[38;2;250;217;83mp[38;2;248;218;91mp[38;2;216;193;85mO[38;2;231;220;122md[38;2;251;237;120mh[38;2;253;229;96mb[38;2;181;162;83mC[38;2;15;9;3m.[38;2;165;150;81mY[38;2;232;207;106mq[38;2;83;73;33m_[38;2;41;36;24mI[38;2;61;52;36mi[38;2;154;144;92mY[38;2;144;126;54mu[38;2;169;142;79mY[38;2;119;89;43mf[38;2;170;147;81mY[38;2;106;94;51mf[38;2;160;157;148mQ[38;2;202;193;180md[38;2;221;204;177mk[38;2;235;219;186mo[38;2;221;205;171mk[38;2;206;190;154mp[38;2;218;203;160mb[38;2;242;225;174mo[38;2;253;231;173m*[38;2;254;224;168m*[38;2;253;220;169mo[38;2;251;225;183m*[38;2;253;245;214m&[38;2;255;252;227mB[38;2;201;191;170mp[38;2;123;110;88mu[38;2;109;99;75mr[38;2;85;78;57m?[38;2;42;40;32ml[38;2;4;4;4m [38;2;0;0;0m    [38;2;7;3;3m [38;2;15;11;9m'[38;2;22;18;15m^[38;2;19;15;12m^[38;2;20;16;13m^[38;2;13;8;6m.[38;2;11;6;5m.[38;2;10;7;6m.[38;2;10;8;7m.[38;2;6;5;4m..[38;2;5;4;3m [38;2;0;0;0m [38;2;0;0;1m [38;2;2;2;1m [38;2;0;0;1m [38;2;25;20;16m\"[38;2;149;134;110mY[38;2;202;181;142mw[38;2;170;148;107mJ[38;2;114;97;76mr[38;2;13;7;3m.[38;2;123;117;72mn[38;2;141;134;72mc[38;2;117;109;64mx[38;2;97;88;53mt[38;2;90;83;51m1[38;2;89;83;49m?[38;2;88;82;51m?[38;2;80;74;43m-[38;2;73;67;36m+[38;2;77;71;40m_[38;2;110;102;55mj[38;2;154;141;76mz[38;2;170;152;75mY[38;2;196;175;81mL[38;2;217;193;88mZ[38;2;211;187;79m0[38;2;216;193;80mO[38;2;231;211;92mw[38;2;189;171;93mQ[38;2;142;130;108mX[38;2;168;164;161mO[38;2;254;253;242m@[38;2;255;251;239m@[38;2;255;247;233mB[38;2;255;248;231mB[38;2;255;249;219m8[38;2;249;235;195mM[38;2;203;186;148mq[38;2;156;139;111mU[38;2;191;176;156mw[38;2;235;228;205m#[38;2;255;249;231mB[38;2;255;247;223m8[38;2;255;240;214m&[38;2;252;236;207mW[38;2;197;181;155mw[38;2;132;116;94mv[38;2;167;152;126mL[38;2;171;155;128mQ[38;2;207;191;164mp[38;2;236;222;191m*[38;2;179;168;139mO[38;2;130;119;98mc[38;2;193;184;163mq[38;2;191;184;157mw[38;2;230;220;191mo[38;2;237;223;199m*[38;2;223;208;180mh[38;2;224;204;164mk[38;2;232;207;160mk[38;2;242;213;158mh[38;2;231;203;144mb[38;2;186;153;117mQ[38;2;149;113;85mc[38;2;177;150;116mL[38;2;104;89;69mj[38;2;91;84;74mf[38;2;49;45;36m![38;2;38;36;28mI[38;2;25;23;19m\"[38;2;8;6;7m.[38;2;0;0;0m                                  [38;2;0;0;0m");
  $display("[38;2;0;0;0m [38;2;1;1;2m [38;2;82;80;56m?[38;2;227;214;126md[38;2;244;219;108md[38;2;249;220;102md[38;2;247;219;92mp[38;2;246;217;83mq[38;2;247;218;85mp[38;2;247;216;85mq[38;2;246;216;84mq[38;2;247;215;87mp[38;2;246;216;87mp[38;2;247;217;86mp[38;2;251;217;88mp[38;2;239;208;93mq[38;2;199;180;89m0[38;2;247;240;153mo[38;2;250;232;119mk[38;2;251;223;105mb[38;2;138;116;69mu[38;2;5;0;0m [38;2;166;151;77mY[38;2;201;176;84mQ[38;2;66;52;27mi[38;2;69;61;46m+[38;2;81;69;41m_[38;2;132;122;74mu[38;2;141;123;54mu[38;2;192;166;79mC[38;2;156;128;45mu[38;2;190;169;83mL[38;2;104;94;52mf[38;2;153;151;145mL[38;2;217;211;197ma[38;2;180;166;138mO[38;2;197;180;146mw[38;2;166;149;121mC[38;2;123;106;90mu[38;2;119;104;85mn[38;2;135;121;93mc[38;2;188;175;138mZ[38;2;223;211;174mh[38;2;233;221;190mo[38;2;239;232;212mM[38;2;230;230;216mM[38;2;178;173;159mm[38;2;134;123;106mz[38;2;113;102;84mx[38;2;116;107;86mn[38;2;135;129;108mX[38;2;139;135;121mY[38;2;88;86;78mf[38;2;64;62;58m_[38;2;50;49;48mi[38;2;44;44;43m![38;2;32;34;30mI[38;2;13;16;13m^[38;2;6;9;6m.[38;2;2;4;4m [38;2;2;3;4m [38;2;4;5;5m [38;2;6;7;7m.[38;2;6;6;7m.[38;2;5;4;5m  [38;2;2;2;3m [38;2;2;2;2m [38;2;1;1;1m [38;2;0;0;0m     [38;2;47;37;29ml[38;2;166;152;121mC[38;2;189;166;126mO[38;2;176;152;127mQ[38;2;19;8;6m'[38;2;136;123;70mu[38;2;239;218;109md[38;2;230;206;97mw[38;2;221;194;92mZ[38;2;203;179;87m0[38;2;187;164;77mC[38;2;180;159;77mJ[38;2;171;150;72mY[38;2;162;139;65mz[38;2;158;135;63mc[38;2;154;131;56mv[38;2;153;130;52mv[38;2;163;138;56mz[38;2;173;149;59mX[38;2;184;161;67mU[38;2;193;170;71mC[38;2;195;171;73mC[38;2;185;166;81mC[38;2;147;136;88mz[38;2;136;131;114mX[38;2;248;246;236mB[38;2;255;252;239m@[38;2;255;249;233mB[38;2;255;239;222m8[38;2;230;211;183ma[38;2;199;182;148mw[38;2;187;173;138mZ[38;2;178;166;140mO[38;2;151;140;125mJ[38;2;155;147;134mC[38;2;240;233;214mW[38;2;253;241;213m&[38;2;248;229;187m#[38;2;250;223;173m*[38;2;246;214;168ma[38;2;187;156;120mQ[38;2;168;145;114mC[38;2;196;179;143mm[38;2;245;231;196mM[38;2;255;246;212m&[38;2;247;234;195mM[38;2;239;228;197m#[38;2;200;192;171mp[38;2;152;143;131mC[38;2;175;165;141mO[38;2;188;175;137mZ[38;2;158;140;113mU[38;2;186;165;135mO[38;2;236;209;166mh[38;2;214;182;136mw[38;2;182;146;100mC[38;2;173;132;84mY[38;2;197;145;88mC[38;2;240;189;114mq[38;2;195;159;99mQ[38;2;103;86;66mf[38;2;168;166;163mZ[38;2;12;12;15m'[38;2;0;0;0m                                     [38;2;0;0;0m");
  $display("[38;2;0;0;0m  [38;2;41;35;26mI[38;2;180;159;86mJ[38;2;209;181;74mQ[38;2;213;184;78m0[38;2;221;193;78mO[38;2;234;207;88mw[38;2;239;211;86mw[38;2;243;213;86mq[38;2;246;216;84mq[38;2;247;217;86mpp[38;2;246;217;84mq[38;2;249;216;84mp[38;2;241;211;89mq[38;2;190;170;81mL[38;2;241;235;149ma[38;2;251;235;120mh[38;2;252;226;107mb[38;2;122;108;65mx[38;2;0;0;0m [38;2;145;130;73mc[38;2;238;220;115md[38;2;112;98;47mf[38;2;64;54;32mi[38;2;90;77;45m?[38;2;102;90;58mf[38;2;149;131;66mc[38;2;228;205;91mw[38;2;213;189;74m0[38;2;187;172;91mL[38;2;60;52;29mi[38;2;136;131;133mU[38;2;255;255;255m$[38;2;216;206;180mk[38;2;220;204;163mb[38;2;232;215;178ma[38;2;146;132;110mY[38;2;53;43;34m![38;2;56;51;45mi[38;2;65;63;54m_[38;2;91;92;85mj[38;2;108;109;104mu[38;2;109;110;107mu[38;2;93;93;91mr[38;2;65;65;61m_[38;2;55;55;51m~[38;2;40;39;37ml[38;2;31;30;28m;[38;2;32;31;28m;[38;2;34;32;29m;[38;2;47;46;43m![38;2;61;62;58m_[38;2;69;71;67m?[38;2;77;81;74m1[38;2;100;107;99mn[38;2;106;110;103mu[38;2;97;101;95mx[38;2;82;85;82mf[38;2;77;79;78mt[38;2;74;76;73m1[38;2;66;66;64m-[38;2;58;58;58m+[38;2;39;39;39ml[38;2;31;31;31m;;[38;2;20;20;20m\"[38;2;19;19;19m\"[38;2;18;18;18m^[38;2;20;20;20m\"[38;2;13;13;13m'[38;2;9;9;9m.[38;2;8;9;10m.[38;2;10;9;9m.[38;2;47;44;36m![38;2;100;88;69mf[38;2;154;140;127mJ[38;2;19;16;13m^[38;2;63;55;30mi[38;2;214;194;103mm[38;2;220;195;84mZ[38;2;217;192;77mO[38;2;209;187;77m0[38;2;198;175;76mL[38;2;188;167;75mC[38;2;179;158;72mU[38;2;164;141;62mz[38;2;169;145;73mY[38;2;163;139;67mz[38;2;150;127;53mv[38;2;155;132;54mv[38;2;177;156;69mU[38;2;187;164;73mJ[38;2;191;165;67mJ[38;2;226;201;97mw[38;2;164;147;87mY[38;2;138;133;118mY[38;2;216;213;200ma[38;2;254;253;238m@[38;2;245;242;225m&[38;2;211;194;172mb[38;2;167;140;111mJ[38;2;193;165;126mO[38;2;222;201;158mb[38;2;242;227;187m*[38;2;255;245;210m&[38;2;255;245;219m8[38;2;177;164;140mO[38;2;202;180;145mw[38;2;253;226;179m*[38;2;232;202;148mb[38;2;197;164;121mO[38;2;179;148;112mC[38;2;201;173;128mZ[38;2;250;223;172m*[38;2;237;209;160mh[38;2;218;193;141mp[38;2;204;176;124mZ[38;2;189;158;103mL[38;2;201;171;117mO[38;2;199;169;117mO[38;2;178;147;110mC[38;2;157;131;89mX[38;2;201;183;132mm[38;2;164;149;118mC[38;2;101;90;74mj[38;2;84;61;47m-[38;2;169;133;87mY[38;2;225;178;111mm[38;2;237;188;117mq[38;2;236;188;113mq[38;2;243;202;130md[38;2;211;183;133mw[38;2;200;187;160mq[38;2;232;230;218mM[38;2;44;44;46m![38;2;0;0;0m                                     [38;2;0;0;0m");
  $display("[38;2;32;32;37mI[38;2;93;91;101mr[38;2;81;73;56m?[38;2;178;158;87mJ[38;2;212;189;89mO[38;2;207;185;79m0[38;2;198;175;69mL[38;2;202;177;74mQ[38;2;200;172;70mL[38;2;205;174;71mL[38;2;218;188;76mO[38;2;231;204;87mw[38;2;242;216;91mp[38;2;247;220;87mp[38;2;244;218;84mq[38;2;247;218;90mp[38;2;207;181;82m0[38;2;214;206;118mq[38;2;255;238;124mh[38;2;255;232;105mk[38;2;152;138;74mz[38;2;7;7;4m.[38;2;51;45;24ml[38;2;225;211;110mq[38;2;189;174;90mQ[38;2;54;42;21ml[38;2;70;61;39m+[38;2;78;71;43m-[38;2;90;81;47m?[38;2;116;106;58mr[38;2;89;80;41m?[38;2;50;43;29ml[38;2;14;11;11m'[38;2;94;90;92mr[38;2;157;157;155m0[38;2;114;112;104mv[38;2;65;60;49m+[38;2;59;54;46m~[38;2;69;67;63m-[38;2;65;64;61m_[38;2;58;56;53m+[38;2;37;36;34mI[38;2;14;15;15m^[38;2;9;9;10m.[38;2;3;3;3m [38;2;0;0;0m  [38;2;1;2;1m [38;2;15;18;17m^[38;2;34;37;35mI[38;2;59;62;58m+[38;2;81;84;79mt[38;2;96;99;94mx[38;2;99;102;95mx[38;2;97;100;91mx[38;2;88;91;83mj[38;2;70;73;65m?[38;2;63;66;59m_[38;2;51;53;49m~[38;2;25;26;25m,[38;2;18;19;19m^[38;2;14;14;14m^[38;2;7;7;7m.[38;2;6;6;6m.[38;2;4;4;4m [38;2;1;1;1m [38;2;3;3;3m [38;2;1;1;1m [38;2;2;2;2m [38;2;3;3;3m [38;2;8;8;8m.[38;2;7;7;7m.[38;2;6;6;6m.[38;2;9;9;9m.[38;2;25;25;25m,[38;2;33;35;36mI[38;2;30;28;29m;[38;2;22;19;18m\"[38;2;5;5;4m [38;2;15;9;5m.[38;2;155;139;75mz[38;2;194;170;76mC[38;2;196;171;72mC[38;2;180;156;62mY[38;2;168;143;61mX[38;2;153;128;55mv[38;2;147;123;56mu[38;2;142;119;55mn[38;2;147;123;60mv[38;2;145;122;55mu[38;2;166;144;72mX[38;2;171;148;72mY[38;2;180;157;75mU[38;2;164;142;56mz[38;2;178;157;70mU[38;2;173;153;85mU[38;2;136;124;99mz[38;2;189;188;180mp[38;2;234;235;222mW[38;2;255;253;241m@[38;2;155;149;134mC[38;2;180;160;132m0[38;2;209;176;128mm[38;2;214;180;125mm[38;2;229;199;145md[38;2;240;215;164ma[38;2;230;206;161mk[38;2;213;191;149mp[38;2;211;192;148mp[38;2;213;190;147mp[38;2;190;164;124m0[38;2;190;162;122m0[38;2;217;188;144mp[38;2;247;223;173mo[38;2;255;233;171m*[38;2;252;222;148ma[38;2;233;190;119mq[38;2;192;140;71mU[38;2;218;160;86mQ[38;2;243;180;104mw[38;2;248;192;111mp[38;2;246;191;111mq[38;2;201;154;98mQ[38;2;102;70;41m?[38;2;58;43;28m![38;2;27;17;10m^[38;2;103;89;70mj[38;2;127;104;67mx[38;2;150;116;71mv[38;2;173;133;85mY[38;2;182;145;94mJ[38;2;189;156;103mL[38;2;219;193;142mp[38;2;238;220;183mo[38;2;240;229;208mM[38;2;202;195;178md[38;2;62;59;57m+[38;2;25;24;28m,[38;2;0;0;0m                                    [38;2;0;0;0m");
  $display("[38;2;40;38;41ml[38;2;110;105;100mn[38;2;120;112;71mn[38;2;167;150;85mU[38;2;154;134;62mc[38;2;158;137;52mc[38;2;180;158;64mU[38;2;192;169;68mC[38;2;196;173;70mC[38;2;205;180;80mQ[38;2;198;172;73mL[38;2;190;165;66mJ[38;2;202;178;68mL[38;2;222;197;75mO[38;2;238;214;89mq[38;2;245;218;89mp[38;2;241;213;95mp[38;2;185;167;70mJ[38;2;240;220;118mb[38;2;255;236;107mk[38;2;197;183;93m0[38;2;20;18;9m^[38;2;0;0;0m [38;2;101;87;51mt[38;2;194;180;106mO[38;2;111;98;64mj[38;2;38;30;25m;[38;2;8;6;6m.[38;2;0;0;0m  [38;2;0;0;1m [38;2;0;0;0m [38;2;5;5;6m.[38;2;3;3;4m [38;2;0;0;0m   [38;2;7;8;9m.[38;2;17;18;19m^[38;2;3;3;3m [38;2;0;0;0m     [38;2;1;2;0m [38;2;10;12;9m'[38;2;44;47;44m![38;2;81;86;82mf[38;2;102;108;101mn[38;2;106;113;105mu[38;2;100;107;99mn[38;2;83;88;80mf[38;2;57;60;54m+[38;2;28;29;27m;[38;2;9;9;9m.[38;2;2;2;2m [38;2;0;0;0m          [38;2;1;1;1m   [38;2;0;0;0m     [38;2;2;2;2m [38;2;9;9;9m.[38;2;11;11;12m'[38;2;1;1;3m [38;2;7;5;6m.[38;2;65;59;38m~[38;2;109;94;54mf[38;2;169;149;76mY[38;2;202;177;84mQ[38;2;199;170;78mL[38;2;189;162;71mJ[38;2;188;163;77mC[38;2;163;138;64mz[38;2;159;135;69mz[38;2;155;133;66mc[38;2;161;143;68mX[38;2;172;153;73mY[38;2;180;157;75mU[38;2;179;157;72mU[38;2;162;146;78mY[38;2;100;85;65mf[38;2;97;88;80mj[38;2;167;164;154mO[38;2;253;251;239m@[38;2;255;252;235m@[38;2;189;180;158mw[38;2;178;161;125mQ[38;2;218;192;144mp[38;2;234;207;160mk[38;2;207;182;141mw[38;2;185;164;126m0[38;2;174;152;115mL[38;2;156;134;100mY[38;2;150;131;103mY[38;2;168;148;118mC[38;2;197;174;139mm[38;2;250;228;176m*[38;2;253;233;177m#[38;2;226;208;156mb[38;2;216;199;149md[38;2;184;160;114mQ[38;2;133;101;60mx[38;2;183;141;90mJ[38;2;217;172;104mO[38;2;207;163;102m0[38;2;167;129;85mX[38;2;181;148;105mC[38;2;166;139;104mU[38;2;164;142;119mJ[38;2;165;152;129mL[38;2;148;139;113mU[38;2;127;115;91mv[38;2;144;132;100mX[38;2;205;189;153mq[38;2;210;190;150mp[38;2;219;197;158md[38;2;220;201;161mb[38;2;222;207;167mk[38;2;228;213;179ma[38;2;233;217;190mo[38;2;235;220;195m*[38;2;191;177;163mw[38;2;112;105;97mn[38;2;61;60;56m+[38;2;4;4;4m [38;2;0;0;0m                                  [38;2;0;0;0m");
  $display("[38;2;37;38;26mI[38;2;174;170;118mQ[38;2;222;216;124mp[38;2;225;211;120mp[38;2;212;196;109mm[38;2;192;173;80mL[38;2;183;164;69mJ[38;2;186;165;71mJ[38;2;173;150;57mX[38;2;170;147;58mX[38;2;180;158;67mU[38;2;176;155;61mY[38;2;185;162;66mU[38;2;190;165;68mJ[38;2;205;177;76mQ[38;2;223;195;79mZ[38;2;245;219;90mp[38;2;224;200;90mm[38;2;198;173;84mQ[38;2;254;238;132ma[38;2;244;232;145ma[38;2;69;65;44m+[38;2;0;0;0m [38;2;30;24;12m\"[38;2;133;113;62mn[38;2;203;181;92m0[38;2;200;183;99mO[38;2;86;79;47m?[38;2;5;4;3m [38;2;0;0;1m [38;2;1;0;4m [38;2;1;1;2m [38;2;0;0;1m [38;2;0;0;0m [38;2;1;1;1m  [38;2;0;0;0m    [38;2;1;1;1m [38;2;0;0;0m  [38;2;1;1;1m  [38;2;1;2;0m [38;2;16;18;15m^[38;2;57;59;55m+[38;2;87;89;84mf[38;2;89;92;86mj[38;2;66;71;65m-[38;2;38;44;38ml[38;2;14;16;13m^[38;2;3;3;3m [38;2;0;0;0m                       [38;2;0;0;1m [38;2;1;1;3m [38;2;2;1;4m [38;2;0;0;2m  [38;2;44;39;25mI[38;2;134;119;67mu[38;2;196;174;89mQ[38;2;228;206;97mw[38;2;236;213;95mq[38;2;233;210;94mq[38;2;203;179;85mQ[38;2;157;135;63mc[38;2;144;126;59mu[38;2;157;139;68mz[38;2;148;127;57mv[38;2;142;126;64mv[38;2;90;81;51m1[38;2;92;83;83mf[38;2;67;61;50m+[38;2;185;179;164mw[38;2;248;239;216m&[38;2;237;226;193m*[38;2;198;184;146mw[38;2;145;129;96mz[38;2;111;91;72mj[38;2;104;86;72mj[38;2;68;54;41m~[38;2;130;117;102mc[38;2;204;192;170md[38;2;206;193;167md[38;2;224;209;182mh[38;2;238;219;184mo[38;2;244;224;178m*[38;2;244;224;174mo[38;2;170;154;121mL[38;2;191;179;164mw[38;2;233;225;218mM[38;2;188;178;165mw[38;2;171;156;133mQ[38;2;226;204;166mk[38;2;232;204;159mk[38;2;236;207;171mh[38;2;182;155;126mQ[38;2;185;160;124m0[38;2;250;228;186m#[38;2;250;232;191mM[38;2;252;241;205mW[38;2;251;246;216m&[38;2;201;194;180md[38;2;107;100;87mx[38;2;206;199;183mb[38;2;255;254;234m@[38;2;255;245;223m8[38;2;254;243;220m8[38;2;254;242;219m8[38;2;255;243;222m8[38;2;255;245;224m8[38;2;255;247;231mB[38;2;249;239;225m&[38;2;121;114;98mv[38;2;100;98;84mr[38;2;32;32;28m;[38;2;0;0;0m                                  [38;2;0;0;0m");
  $display("[38;2;33;33;23m;[38;2;118;112;73mn[38;2;146;130;75mc[38;2;158;137;78mX[38;2;186;167;103mQ[38;2;206;190;115mm[38;2;214;202;115mw[38;2;230;220;125md[38;2;238;225;125mb[38;2;226;211;111mq[38;2;200;185;88m0[38;2;180;163;71mJ[38;2;172;152;61mY[38;2;166;143;49mz[38;2;177;151;63mY[38;2;188;160;68mJ[38;2;201;176;68mL[38;2;228;202;92mw[38;2;194;171;82mL[38;2;221;210;127mp[38;2;237;234;161ma[38;2;136;135;99mz[38;2;9;4;2m.[38;2;136;126;69mv[38;2;242;221;105md[38;2;251;223;92md[38;2;252;228;92md[38;2;251;237;128mh[38;2;181;176;120m0[38;2;61;61;47m+[38;2;0;0;0m           [38;2;1;0;0m [38;2;0;0;0m  [38;2;1;1;1m  [38;2;5;6;5m.[38;2;30;31;29m;[38;2;75;76;74m1[38;2;80;81;78mt[38;2;15;17;16m^[38;2;0;1;1m [38;2;1;2;2m [38;2;1;1;1m  [38;2;0;0;0m                  [38;2;1;1;1m    [38;2;0;0;1m [38;2;2;2;3m [38;2;1;1;3m  [38;2;0;0;3m [38;2;1;0;3m [38;2;8;4;7m.[38;2;24;19;11m^[38;2;63;54;30mi[38;2;119;108;56mr[38;2;189;178;90mQ[38;2;198;183;95m0[38;2;145;129;60mv[38;2;131;115;59mn[38;2;116;101;42mf[38;2;117;101;50mj[38;2;96;83;55mt[38;2;100;90;81mj[38;2;75;66;55m-[38;2;117;105;82mn[38;2;157;139;110mU[38;2;177;157;120mQ[38;2;156;134;96mY[38;2;168;146;111mJ[38;2;145;122;95mz[38;2;122;100;77mx[38;2;118;101;78mx[38;2;195;182;157mw[38;2;253;240;212m&[38;2;255;244;216m8[38;2;255;242;212m&[38;2;255;237;205mW[38;2;255;230;190mM[38;2;255;232;172m*[38;2;232;214;161mh[38;2;149;139;113mU[38;2;255;250;238m@[38;2;254;252;240m@[38;2;255;255;245m@[38;2;208;205;194mh[38;2;211;204;191mh[38;2;252;245;223m8[38;2;251;243;215m&[38;2;230;221;195m*[38;2;197;188;169mp[38;2;253;244;227m8[38;2;254;245;228m8[38;2;255;250;232mB[38;2;255;251;228mB[38;2;254;246;221m8[38;2;134;123;101mz[38;2;147;128;109mY[38;2;185;159;129m0[38;2;193;162;117m0[38;2;209;176;123mZ[38;2;216;182;131mw[38;2;224;196;153md[38;2;223;199;163mb[38;2;230;213;182ma[38;2;207;194;167md[38;2;163;154;128mL[38;2;119;110;88mn[38;2;126;118;103mc[38;2;88;87;80mf[38;2;1;1;0m [38;2;0;0;0m                                [38;2;0;0;0m");
  $display("[38;2;67;62;35m~[38;2;227;215;124md[38;2;242;225;114mb[38;2;240;223;111md[38;2;232;217;112mp[38;2;205;194;109mZ[38;2;159;152;90mU[38;2;130;125;79mv[38;2;123;117;72mn[38;2;148;141;86mX[38;2;194;184;112mO[38;2;228;219;122md[38;2;240;229;118mb[38;2;230;214;106mp[38;2;211;191;85mO[38;2;203;181;78mQ[38;2;194;171;67mC[38;2;188;164;59mU[38;2;198;176;78mL[38;2;193;182;95m0[38;2;242;240;159mo[38;2;229;230;166ma[38;2;70;64;44m+[38;2;98;89;42m1[38;2;216;194;91mZ[38;2;250;220;97md[38;2;251;224;88mp[38;2;255;234;108mk[38;2;255;247;139mo[38;2;242;235;158mo[38;2;158;152;109mJ[38;2;76;73;53m-[38;2;59;55;42m~[38;2;60;58;45m~[38;2;57;54;42m~[38;2;34;30;23m;[38;2;15;12;10m'[38;2;5;4;2m [38;2;0;0;0m        [38;2;7;7;7m.[38;2;22;22;22m\"[38;2;39;39;39mll[38;2;10;10;10m'[38;2;1;1;1m  [38;2;0;0;0m                   [38;2;1;1;1m   [38;2;0;0;0m    [38;2;1;1;1m [38;2;1;1;2m [38;2;0;0;1m [38;2;2;1;1m [38;2;9;9;9m.[38;2;14;14;14m^[38;2;9;10;11m'[38;2;0;0;0m [38;2;18;15;14m^[38;2;67;62;41m+[38;2;100;92;56mt[38;2;94;81;39m?[38;2;118;105;52mj[38;2;115;102;67mr[38;2;157;146;129mC[38;2;109;98;81mx[38;2;126;113;91mv[38;2;158;139;107mU[38;2;163;137;92mY[38;2;179;152;101mC[38;2;206;181;125mm[38;2;220;198;145mp[38;2;173;151;110mC[38;2;168;146;108mJ[38;2;209;188;149mq[38;2;229;210;171mh[38;2;243;227;186m*[38;2;252;235;192mM[38;2;253;233;188mM[38;2;252;227;180m*[38;2;253;227;178m*[38;2;234;212;159mk[38;2;198;184;142mw[38;2;148;140;119mU[38;2;204;198;183mb[38;2;250;245;231m8[38;2;255;248;233mB[38;2;255;248;231mB[38;2;231;223;203m*[38;2;230;223;199m*[38;2;225;219;191mo[38;2;220;214;191ma[38;2;239;232;209mM[38;2;244;233;212mW[38;2;231;217;193mo[38;2;212;189;157mp[38;2;204;174;132mm[38;2;215;180;127mw[38;2;197;167;116mO[38;2;143;114;81mv[38;2;164;134;99mY[38;2;186;151;103mC[38;2;185;149;98mC[38;2;187;152;106mL[38;2;184;156;119mQ[38;2;174;155;124mQ[38;2;183;168;139mO[38;2;178;166;140mO[38;2;134;124;101mz[38;2;199;188;166mp[38;2;221;209;190ma[38;2;155;150;137mL[38;2;23;22;22m\"[38;2;5;6;8m.[38;2;0;1;3m [38;2;0;0;0m                              [38;2;0;0;0m");
  $display("[38;2;71;66;35m+[38;2;240;224;126mb[38;2;253;234;113mk[38;2;255;235;113mk[38;2;255;236;109mk[38;2;253;238;112mk[38;2;253;241;124ma[38;2;249;238;137ma[38;2;208;198;124mw[38;2;142;134;87mz[38;2;87;81;51m?[38;2;64;58;36m~[38;2;74;66;38m+[38;2;129;119;69mn[38;2;195;183;103mO[38;2;225;212;114mp[38;2;242;228;119mb[38;2;239;223;103md[38;2;230;213;99mq[38;2;179;165;76mJ[38;2;234;224;142mk[38;2;255;251;169mM[38;2;180;174;127mO[38;2;50;41;25ml[38;2;94;75;45m?[38;2;167;144;75mY[38;2;209;188;79m0[38;2;238;216;93mq[38;2;249;229;96md[38;2;251;232;105mb[38;2;255;241;133ma[38;2;255;240;153m*[38;2;252;237;161m*[38;2;253;240;170m#[38;2;250;241;172m#[38;2;236;229;162ma[38;2;214;208;147md[38;2;195;189;129mm[38;2;168;165;102mC[38;2;140;136;81mz[38;2;82;77;46m-[38;2;24;20;14m\"[38;2;10;9;12m'[38;2;18;19;19m^[38;2;15;15;15m^[38;2;10;10;10m'[38;2;2;2;2m [38;2;0;0;0m                       [38;2;1;1;1m     [38;2;0;0;0m [38;2;1;1;1m       [38;2;0;0;0m [38;2;1;1;1m [38;2;4;4;5m [38;2;3;4;3m [38;2;0;0;3m [38;2;0;0;0m [38;2;21;17;15m^[38;2;37;30;21m;[38;2;103;95;71mj[38;2;180;170;151mZ[38;2;189;179;163mw[38;2;139;127;99mz[38;2;172;153;117mL[38;2;180;153;108mL[38;2;195;166;110m0[38;2;217;187;127mw[38;2;180;152;102mC[38;2;151;125;89mz[38;2;168;145;110mJ[38;2;181;159;119mQ[38;2;184;162;121mQ[38;2;186;166;122m0[38;2;206;187;137mw[38;2;236;214;163mh[38;2;249;224;172m*[38;2;244;221;170mo[38;2;196;182;142mm[38;2;127;117;102mc[38;2;198;193;184md[38;2;233;228;211mM[38;2;193;182;161mw[38;2;162;146;122mC[38;2;172;151;121mL[38;2;155;133;99mY[38;2;159;138;103mU[38;2;148;127;97mX[38;2;134;111;85mv[38;2;149;127;99mX[38;2;146;124;94mz[38;2;153;128;100mX[38;2;177;151;121mL[38;2;200;176;144mm[38;2;229;207;174mh[38;2;239;219;185mo[38;2;225;213;175mh[38;2;141;128;101mz[38;2;168;153;127mL[38;2;241;222;186m*[38;2;240;216;182mo[38;2;244;221;190m*[38;2;248;228;194m#[38;2;253;234;199mM[38;2;255;240;205mW[38;2;255;244;211m&[38;2;184;173;151mZ[38;2;138;125;110mX[38;2;238;225;202m#[38;2;228;219;192mo[38;2;194;188;165mq[38;2;150;145;128mJ[38;2;181;177;163mm[38;2;166;162;147m0[38;2;161;159;145mQ[38;2;70;69;65m-[38;2;2;2;4m [38;2;0;0;0m                          [38;2;0;0;0m");
  $display("[38;2;72;67;34m+[38;2;238;223;122mb[38;2;253;234;111mk[38;2;254;233;115mk[38;2;254;233;117mk[38;2;252;234;113mk[38;2;250;235;115mk[38;2;251;237;121mh[38;2;255;243;138mo[38;2;255;248;153m*[38;2;255;241;150m*[38;2;227;210;125mp[38;2;170;157;83mU[38;2;107;96;50mf[38;2;75;63;44m_[38;2;68;54;36m~[38;2;148;132;82mz[38;2;194;179;96m0[38;2;214;200;112mw[38;2;209;194;114mm[38;2;226;214;133md[38;2;255;248;162m#[38;2;250;246;167m#[38;2;129;122;84mv[38;2;101;91;70mj[38;2;103;92;64mf[38;2;107;95;55mf[38;2;133;119;51mn[38;2;205;185;77mQ[38;2;247;222;94mp[38;2;252;228;101mb[38;2;254;231;115mk[38;2;255;236;132ma[38;2;255;237;142mo[38;2;255;241;150m*[38;2;255;246;160m#[38;2;255;248;166m#[38;2;255;251;167mM[38;2;255;252;156m#[38;2;255;245;136mo[38;2;247;235;124mh[38;2;210;201;107mm[38;2;142;141;88mz[38;2;103;106;91mx[38;2;109;110;108mu[38;2;138;138;133mU[38;2;147;147;145mC[38;2;152;152;150mQ[38;2;151;153;149mQ[38;2;153;155;150mQ[38;2;142;144;141mC[38;2;127;129;126mX[38;2;109;110;108mu[38;2;94;94;92mr[38;2;71;71;70m?[38;2;50;50;48mi[38;2;30;30;28m;[38;2;15;15;15m^[38;2;5;5;5m.[38;2;1;1;1m [38;2;0;0;0m   [38;2;1;1;1m    [38;2;0;0;0m         [38;2;1;1;1m   [38;2;0;0;0m        [38;2;1;2;1m [38;2;1;1;3m [38;2;0;0;1m [38;2;0;0;0m [38;2;87;85;82mf[38;2;212;202;194mh[38;2;171;156;138mQ[38;2;177;158;120mQ[38;2;185;158;110mQ[38;2;187;156;97mC[38;2;184;157;108mL[38;2;155;130;94mX[38;2;152;130;97mX[38;2;171;150;114mC[38;2;179;159;114mL[38;2;180;161;117mQ[38;2;179;160;117mQ[38;2;188;170;125mO[38;2;203;183;136mw[38;2;190;166;121m0[38;2;177;151;110mC[38;2;193;172;135mZ[38;2;203;190;164mp[38;2;238;225;200m#[38;2;246;231;195mM[38;2;242;222;173mo[38;2;245;219;166ma[38;2;233;205;153mk[38;2;210;180;135mw[38;2;191;160;124m0[38;2;178;148;114mC[38;2;178;150;117mL[38;2;192;164;127mO[38;2;217;190;149mp[38;2;238;211;167mh[38;2;249;222;178m*[38;2;255;230;186m#[38;2;255;232;187mM[38;2;253;230;183m#[38;2;248;228;181m*[38;2;247;230;186m#[38;2;160;144;110mJ[38;2;118;96;61mj[38;2;225;198;149md[38;2;241;209;155mk[38;2;232;200;143md[38;2;226;193;138mp[38;2;229;196;145md[38;2;230;200;147mb[38;2;237;213;160mh[38;2;215;192;154mp[38;2;129;105;74mn[38;2;239;215;171ma[38;2;243;221;168ma[38;2;230;209;155mk[38;2;175;153;104mC[38;2;246;222;179m*[38;2;255;237;192mM[38;2;255;241;202mW[38;2;201;189;169mp[38;2;26;24;22m,[38;2;0;0;0m                          [38;2;0;0;0m");
  $display("[38;2;74;68;35m+[38;2;240;224;120mb[38;2;254;235;108mk[38;2;254;235;110mk[38;2;255;235;112mk[38;2;252;235;111mkk[38;2;254;235;115mk[38;2;252;235;128mh[38;2;254;237;144mo[38;2;255;240;151m*[38;2;255;243;144mo[38;2;255;242;131ma[38;2;247;230;115mk[38;2;218;198;93mZ[38;2;155;134;69mz[38;2;113;92;51mf[38;2;155;139;83mX[38;2;190;171;97mQ[38;2;195;175;99m0[38;2;191;177;110m0[38;2;214;205;141mp[38;2;245;239;170m*[38;2;216;207;156mb[38;2;102;94;65mj[38;2;203;201;148mp[38;2;169;166;114mL[38;2;121;112;77mn[38;2;103;84;46m1[38;2;162;139;68mz[38;2;218;196;88mZ[38;2;245;225;92mp[38;2;250;232;102mb[38;2;253;236;119mh[38;2;254;237;125mh[38;2;253;237;139ma[38;2;254;238;151mo[38;2;255;241;159m*[38;2;253;244;153m*[38;2;254;243;145mo[38;2;253;238;122mh[38;2;255;237;105mk[38;2;252;237;118mh[38;2;186;175;95mQ[38;2;51;48;27m![38;2;13;13;14m'[38;2;37;38;38ml[38;2;47;47;46mi[38;2;50;51;48mi[38;2;54;54;53m~[38;2;59;59;58m+[38;2;68;68;66m-[38;2;77;77;76m1[38;2;88;88;87mj[38;2;94;95;94mr[38;2;97;97;96mx[38;2;112;112;111mv[38;2;118;119;117mc[38;2;103;105;102mn[38;2;102;104;100mn[38;2;113;115;111mv[38;2;84;85;81mf[38;2;24;25;23m,[38;2;3;3;2m [38;2;0;0;0m  [38;2;1;1;1m [38;2;0;0;0m  [38;2;1;1;1m [38;2;0;0;0m     [38;2;1;1;1m  [38;2;0;0;0m [38;2;6;6;6m.[38;2;9;9;9m.[38;2;11;11;11m'[38;2;14;14;14m^[38;2;18;18;18m^[38;2;12;12;12m'[38;2;8;8;8m.[38;2;13;13;13m'[38;2;11;11;12m'[38;2;7;7;7m.[38;2;4;4;4m [38;2;0;0;0m [38;2;38;40;37ml[38;2;151;151;142mL[38;2;185;176;157mm[38;2;196;179;149mw[38;2;197;172;129mZ[38;2;196;169;121mO[38;2;180;157;111mL[38;2;159;142;113mJ[38;2;192;178;161mw[38;2;221;208;185mh[38;2;221;205;171mk[38;2;221;203;162mb[38;2;190;171;132mO[38;2;192;174;134mZ[38;2;184;165;128m0[38;2;160;140;104mU[38;2;152;128;90mz[38;2;180;153;111mL[38;2;214;184;138mw[38;2;212;184;133mw[38;2;217;188;135mq[38;2;242;210;155mh[38;2;250;219;162ma[38;2;246;217;157ma[38;2;248;216;157ma[38;2;250;218;162ma[38;2;252;220;164mo[38;2;249;218;161ma[38;2;247;217;159ma[38;2;254;222;167mo[38;2;255;222;169m*[38;2;249;216;164ma[38;2;236;205;155mk[38;2;221;194;144mp[38;2;207;180;127mm[38;2;215;181;127mw[38;2;216;183;126mw[38;2;200;170;115mO[38;2;182;155;107mL[38;2;161;130;80mz[38;2;187;145;85mJ[38;2;213;165;95m0[38;2;213;166;94m0[38;2;210;166;94m0[38;2;215;173;103mO[38;2;215;178;109mZ[38;2;204;170;114mO[38;2;154;120;81mc[38;2;169;136;94mU[38;2;216;184;127mw[38;2;206;174;108mO[38;2;207;174;108mO[38;2;214;178;119mm[38;2;208;170;121mZ[38;2;200;168;126mO[38;2;177;157;124mQ[38;2;92;87;72mf[38;2;8;8;8m.[38;2;0;0;0m                          [38;2;0;0;0m");
  $display("[38;2;77;72;35m_[38;2;241;225;116mb[38;2;254;235;102mk[38;2;254;235;107mk[38;2;255;234;112mk[38;2;254;234;113mk[38;2;254;234;110mk[38;2;252;235;109mk[38;2;252;235;116mk[38;2;254;235;129ma[38;2;255;237;143mo[38;2;254;239;151mo[38;2;255;239;148mo[38;2;255;239;131ma[38;2;249;229;105mb[38;2;246;222;97md[38;2;216;193;91mZ[38;2;150;128;67mc[38;2;155;134;75mz[38;2;203;179;91m0[38;2;225;202;101mw[38;2;201;181;91m0[38;2;179;167;94mC[38;2;174;167;114mQ[38;2;94;89;56mt[38;2;216;214;139md[38;2;253;247;159m*[38;2;240;228;160ma[38;2;190;177;126mO[38;2;128;113;77mu[38;2;117;100;53mj[38;2;168;148;71mY[38;2;211;189;83mO[38;2;235;215;91mq[38;2;247;227;101md[38;2;252;232;114mk[38;2;255;234;130ma[38;2;255;236;140ma[38;2;254;238;142mo[38;2;254;239;141mo[38;2;254;240;139mo[38;2;253;234;127mh[38;2;250;231;105mb[38;2;255;237;103mk[38;2;226;210;106mq[38;2;93;85;43m?[38;2;0;0;0m           [38;2;3;4;3m [38;2;9;10;9m.[38;2;20;21;19m\"[38;2;35;36;34mI[38;2;69;70;66m-[38;2;77;77;73m1[38;2;62;63;60m_[38;2;35;35;35mI[38;2;13;13;13m'[38;2;3;3;3m [38;2;0;0;0m       [38;2;1;1;1m [38;2;1;1;2m [38;2;6;6;6m.[38;2;18;18;18m^[38;2;30;30;30m;[38;2;31;31;31m;[38;2;33;33;33mI[38;2;28;28;28m;[38;2;17;17;17m^[38;2;11;11;11m''[38;2;12;12;12m'[38;2;9;9;9m.[38;2;4;4;4m [38;2;0;0;0m [38;2;0;0;1m [38;2;103;101;96mx[38;2;207;202;185mk[38;2;222;210;177mh[38;2;211;192;148mp[38;2;214;190;138mq[38;2;213;193;142mq[38;2;183;167;134mO[38;2;231;221;198m*[38;2;255;247;225m8[38;2;255;242;216m&[38;2;255;241;208m&[38;2;249;233;199mM[38;2;191;174;144mZ[38;2;147;129;105mX[38;2;143;124;97mz[38;2;173;153;117mL[38;2;192;170;127mO[38;2;196;170;123mO[38;2;185;150;98mC[38;2;172;135;74mX[38;2;182;149;87mJ[38;2;215;185;134mw[38;2;199;171;132mZ[38;2;216;191;155mp[38;2;220;198;162mb[38;2;222;201;168mk[38;2;216;200;168mb[38;2;209;195;167md[38;2;195;180;152mw[38;2;214;196;166mb[38;2;225;204;169mk[38;2;203;174;130mZ[38;2;180;142;89mU[38;2;199;152;96mL[38;2;216;164;99m0[38;2;225;173;100mZ[38;2;228;180;104mm[38;2;201;156;96mQ[38;2;133;99;54mr[38;2;148;116;75mv[38;2;163;126;81mz[38;2;191;151;98mC[38;2;211;172;114mZ[38;2;218;181;118mm[38;2;220;181;118mm[38;2;216;178;120mm[38;2;199;164;117mO[38;2;169;137;104mU[38;2;128;101;75mn[38;2;167;142;110mJ[38;2;202;172;133mZ[38;2;189;158;115mQ[38;2;159;133;97mY[38;2;113;93;69mj[38;2;87;76;61m1[38;2;45;40;33ml[38;2;4;4;4m [38;2;0;0;1m [38;2;0;0;0m                          [38;2;0;0;0m");
  $display("[38;2;73;68;31m+[38;2;236;220;109md[38;2;252;231;94mb[38;2;254;231;98mb[38;2;254;232;106mk[38;2;254;233;110mk[38;2;254;234;109mk[38;2;254;234;107mk[38;2;254;233;112mk[38;2;253;233;121mh[38;2;253;235;133ma[38;2;254;238;146mo[38;2;254;239;150mo[38;2;254;241;142mo[38;2;253;237;128ma[38;2;246;224;102md[38;2;244;220;94mp[38;2;215;194;94mZ[38;2;136;112;60mn[38;2;183;154;92mC[38;2;189;161;75mJ[38;2;230;203;92mw[38;2;244;222;96mp[38;2;231;212;97mq[38;2;239;222;114md[38;2;250;236;125mh[38;2;249;236;126mh[38;2;252;239;137ma[38;2;255;247;153m*[38;2;244;235;160mo[38;2;187;177;121mO[38;2;150;133;85mz[38;2;148;129;72mc[38;2;150;132;57mv[38;2;187;168;70mJ[38;2;237;215;96mq[38;2;249;229;105mb[38;2;252;234;118mk[38;2;254;235;129ma[38;2;255;236;135ma[38;2;254;237;141ma[38;2;255;237;139ma[38;2;253;234;121mh[38;2;248;229;100mb[38;2;249;229;94md[38;2;242;228;104md[38;2;135;126;66mu[38;2;11;9;5m.[38;2;0;0;2m [38;2;1;1;3m [38;2;0;0;3m [38;2;1;1;4m [38;2;0;0;2m [38;2;0;0;0m          [38;2;10;10;10m'[38;2;28;28;28m;[38;2;41;41;41ml[38;2;48;48;48mi[38;2;41;41;41ml[38;2;40;40;40mll[38;2;29;29;29m;[38;2;20;20;20m\"[38;2;24;24;24m,[38;2;19;19;18m^[38;2;17;17;16m^[38;2;24;24;23m,[38;2;32;32;31m;[38;2;31;31;31m;[38;2;26;26;26m,[38;2;14;14;14m^[38;2;7;7;7m.[38;2;2;2;2m [38;2;0;0;0m [38;2;1;1;1m [38;2;0;0;0m [38;2;1;1;1m [38;2;0;0;0m  [38;2;2;1;2m [38;2;88;84;82mf[38;2;170;162;149mO[38;2;218;209;180mh[38;2;231;215;176ma[38;2;235;214;169ma[38;2;237;213;166mh[38;2;201;183;140mw[38;2;238;225;193m*[38;2;255;244;215m8[38;2;251;239;211mW[38;2;254;239;209m&[38;2;255;240;204mW[38;2;211;195;159md[38;2;155;138;103mY[38;2;179;160;124mQ[38;2;207;186;144mq[38;2;202;180;135mm[38;2;201;177;135mm[38;2;198;174;132mZ[38;2;187;163;118m0[38;2;174;150;105mC[38;2;141;120;83mv[38;2;173;155;132mQ[38;2;213;200;184mk[38;2;247;238;226m&[38;2;249;244;232m8[38;2;249;247;237mB[38;2;252;251;241m@[38;2;255;255;247m$$[38;2;223;220;216m*[38;2;163;155;151m0[38;2;148;133;114mY[38;2;175;149;111mC[38;2;200;167;120mO[38;2;202;167;120mO[38;2;198;170;122mO[38;2;172;146;106mJ[38;2;185;160;134m0[38;2;213;194;172mb[38;2;243;225;197m#[38;2;220;202;169mk[38;2;170;150;116mC[38;2;192;169;128mO[38;2;226;199;153mb[38;2;224;191;144mp[38;2;224;191;145mp[38;2;230;202;156mb[38;2;244;222;180m*[38;2;208;191;159mp[38;2;149;132;103mY[38;2;225;204;163mk[38;2;237;216;170ma[38;2;202;188;153mq[38;2;78;74;59m?[38;2;10;12;13m'[38;2;0;0;0m                             [38;2;0;0;0m");
  $display("[38;2;72;66;30m+[38;2;235;217;104mp[38;2;254;228;88md[38;2;254;229;87md[38;2;254;229;94mb[38;2;254;231;98mb[38;2;253;233;103mb[38;2;254;235;104mk[38;2;254;233;109mk[38;2;254;232;114mk[38;2;254;234;122mh[38;2;254;235;131ma[38;2;254;237;139ma[38;2;253;240;148mo[38;2;254;241;143mo[38;2;253;237;125mh[38;2;242;223;98mp[38;2;247;221;95mp[38;2;204;175;87mQ[38;2;136;109;57mx[38;2;213;185;101mZ[38;2;190;159;75mJ[38;2;200;170;83mQ[38;2;241;216;96mp[38;2;245;222;89mp[38;2;246;226;102md[38;2;252;233;115mk[38;2;254;235;122mh[38;2;252;236;125mh[38;2;253;239;138ma[38;2;254;247;158m*[38;2;227;217;150mk[38;2;180;168;101mL[38;2;180;163;89mC[38;2;149;126;64mv[38;2;149;126;58mv[38;2;207;188;80m0[38;2;241;227;94mp[38;2;250;233;103mb[38;2;254;234;117mk[38;2;254;236;129ma[38;2;253;237;136ma[38;2;255;236;135ma[38;2;253;235;126mh[38;2;249;228;104mb[38;2;248;221;91mp[38;2;249;225;101md[38;2;161;146;79mY[38;2;22;17;10m^[38;2;0;0;0m [38;2;2;1;3m [38;2;1;1;2m [38;2;0;0;1m [38;2;0;0;0m             [38;2;5;5;5m.[38;2;12;12;12m'[38;2;21;21;21m\"[38;2;23;23;23m,[38;2;18;18;18m^[38;2;21;21;21m\"[38;2;19;19;19m\"[38;2;13;13;11m'[38;2;12;13;11m'[38;2;11;11;9m'[38;2;7;7;6m.[38;2;4;4;4m [38;2;1;1;1m [38;2;0;0;0m   [38;2;1;1;1m  [38;2;2;2;2m  [38;2;1;1;1m [38;2;0;0;0m [38;2;68;64;60m-[38;2;189;183;164mw[38;2;231;223;188mo[38;2;241;231;189m#[38;2;250;233;191mM[38;2;244;225;184m*[38;2;197;179;141mm[38;2;235;220;187mo[38;2;255;240;210m&[38;2;251;236;205mW[38;2;252;239;206mW[38;2;249;233;198mM[38;2;208;194;154mp[38;2;205;188;145mq[38;2;230;213;168mh[38;2;238;220;173ma[38;2;240;219;170ma[38;2;243;220;170mo[38;2;228;204;157mb[38;2;186;164;118m0[38;2;175;155;114mL[38;2;133;115;86mv[38;2;175;159;139m0[38;2;250;235;214mW[38;2;255;241;221m8[38;2;251;242;224m8[38;2;254;248;234mB[38;2;253;250;239m@[38;2;254;250;240m@[38;2;255;252;241m@[38;2;249;248;236mB[38;2;142;140;132mJ[38;2;205;202;193mk[38;2;227;222;209m*[38;2;176;168;142mO[38;2;238;228;193m*[38;2;246;233;199mM[38;2;249;237;204mW[38;2;213;199;173mb[38;2;225;212;191ma[38;2;255;247;225m8[38;2;255;249;225mB[38;2;255;255;234m@[38;2;212;206;187mk[38;2;216;208;184mh[38;2;252;239;215m&[38;2;253;238;214m&[38;2;253;241;219m&[38;2;254;245;224m8[38;2;254;249;229mB[38;2;255;254;238m@[38;2;223;218;202mo[38;2;226;219;202m*[38;2;255;252;235m@[38;2;235;226;208m#[38;2;117;109;91mn[38;2;51;45;38m![38;2;6;5;5m.[38;2;0;0;0m                            [38;2;0;0;0m");
  $display("[38;2;66;62;29m~[38;2;231;212;104mq[38;2;255;224;87md[38;2;255;226;86md[38;2;255;229;86md[38;2;254;229;89md[38;2;253;231;96mb[38;2;254;232;101mb[38;2;255;232;106mk[38;2;254;232;108mk[38;2;254;234;114mk[38;2;255;234;120mh[38;2;254;237;128ma[38;2;254;241;147mo[38;2;253;242;153m*[38;2;254;244;141mo[38;2;252;235;120mh[38;2;247;216;94mp[38;2;252;224;96md[38;2;181;161;77mJ[38;2;142;117;60mu[38;2;229;200;106mw[38;2;194;166;80mC[38;2;176;149;72mY[38;2;228;207;93mw[38;2;240;217;91mq[38;2;245;219;98mp[38;2;252;230;115mk[38;2;254;233;120mh[38;2;252;234;124mh[38;2;251;238;131ma[38;2;253;244;151m*[38;2;245;235;159mo[38;2;191;176;106m0[38;2;196;178;97m0[38;2;184;163;88mC[38;2;134;108;50mx[38;2;193;177;80mL[38;2;244;230;96md[38;2;247;228;96md[38;2;253;233;109mk[38;2;254;236;125mh[38;2;255;235;135ma[38;2;254;235;132ma[38;2;255;236;121mh[38;2;251;227;102mb[38;2;246;220;85mp[38;2;251;222;101md[38;2;177;155;86mJ[38;2;28;21;11m\"[38;2;0;0;0m [38;2;1;1;1m  [38;2;0;0;0m           [38;2;1;1;1m [38;2;0;0;0m                   [38;2;1;1;1m [38;2;2;2;2m [38;2;0;0;0m [38;2;39;38;36ml[38;2;166;161;145m0[38;2;234;228;197m*[38;2;246;236;195mM[38;2;250;235;193mM[38;2;244;228;188m#[38;2;194;178;142mm[38;2;229;214;181ma[38;2;255;238;208mW[38;2;253;236;206mW[38;2;255;238;208mW[38;2;239;223;190m*[38;2;196;180;147mw[38;2;224;207;172mk[38;2;255;238;197mW[38;2;255;239;195mW[38;2;255;238;192mM[38;2;255;234;184mM[38;2;245;223;174mo[38;2;238;212;167mh[38;2;180;154;111mL[38;2;145;122;82mc[38;2;170;148;111mC[38;2;219;199;165mb[38;2;231;214;183ma[38;2;236;223;197m*[38;2;250;241;225m8[38;2;255;248;238m@[38;2;255;249;239m@[38;2;254;250;239m@[38;2;253;249;238mB[38;2;253;250;240m@[38;2;209;208;196mh[38;2;185;184;170mq[38;2;251;246;232mB[38;2;221;214;195ma[38;2;190;183;168mq[38;2;200;190;177md[38;2;200;191;171mp[38;2;212;202;181mk[38;2;249;240;217m&[38;2;254;246;220m8[38;2;248;241;214m&[38;2;239;229;207mM[38;2;246;233;212mW[38;2;254;243;219m8[38;2;253;241;221m8[38;2;253;241;223m8[38;2;252;242;224m8[38;2;250;244;225m8[38;2;250;245;226m8[38;2;247;238;219m&[38;2;253;243;216m&[38;2;248;241;216m&[38;2;201;195;181mb[38;2;154;148;133mC[38;2;211;198;175mb[38;2;131;119;99mc[38;2;15;14;14m^[38;2;0;0;0m                            [38;2;0;0;0m");
  $display("[38;2;67;60;29m~[38;2;232;210;104mq[38;2;252;220;86mp[38;2;252;221;85mp[38;2;252;224;83mp[38;2;252;224;84mp[38;2;252;226;90md[38;2;255;229;96mb[38;2;255;231;101mb[38;2;254;232;105mk[38;2;253;233;111mk[38;2;254;233;117mk[38;2;252;234;122mh[38;2;250;237;137ma[38;2;253;242;153m*[38;2;254;243;157m*[38;2;255;241;145mo[38;2;248;225;110mb[38;2;242;217;89mq[38;2;245;223;102md[38;2;177;150;69mY[38;2;178;148;72mY[38;2;235;212;105mp[38;2;206;181;90m0[38;2;167;140;66mX[38;2;225;199;93mm[38;2;247;217;93mp[38;2;246;218;89mp[38;2;252;226;105mb[38;2;254;233;120mh[38;2;251;235;123mh[38;2;248;235;126mh[38;2;253;242;142mo[38;2;251;243;163m*[38;2;195;181;114mO[38;2;195;174;87mQ[38;2;210;190;95mZ[38;2;129;106;47mr[38;2;181;160;76mJ[38;2;245;226;99md[38;2;246;225;92mp[38;2;251;229;105mb[38;2;254;233;120mh[38;2;254;235;125mh[38;2;254;236;125mh[38;2;253;237;116mh[38;2;248;228;99md[38;2;243;218;83mq[38;2;250;220;100md[38;2;183;161;90mC[38;2;32;26;14m,[38;2;0;0;0m [38;2;1;1;3m [38;2;0;0;0m                             [38;2;1;1;1m [38;2;0;0;0m   [38;2;18;18;18m^[38;2;130;127;118mX[38;2;220;213;188ma[38;2;248;238;203mW[38;2;249;236;200mM[38;2;251;235;201mW[38;2;215;198;165mb[38;2;232;216;183ma[38;2;255;239;207mW[38;2;252;236;204mW[38;2;254;237;205mW[38;2;227;211;178mh[38;2;206;191;157mp[38;2;237;223;189m*[38;2;254;238;203mW[38;2;249;235;194mM[38;2;244;229;187m#[38;2;239;221;178mo[38;2;222;202;156mb[38;2;206;181;140mw[38;2;179;151;113mL[38;2;137;107;65mn[38;2;154;119;71mv[38;2;167;131;80mX[38;2;174;144;94mU[38;2;206;184;141mw[38;2;240;230;201m#[38;2;254;249;235mB[38;2;253;249;240m@[38;2;253;251;238m@[38;2;253;250;235mB[38;2;254;249;236mB[38;2;254;248;238mB[38;2;255;251;241m@[38;2;204;194;179mb[38;2;179;158;132m0[38;2;213;191;150mp[38;2;204;183;140mw[38;2;199;177;139mm[38;2;209;187;150mq[38;2;218;195;163mb[38;2;209;184;154mq[38;2;204;182;142mw[38;2;220;200;156mb[38;2;162;143;112mJ[38;2;112;94;76mr[38;2;159;146;121mC[38;2;197;182;148mw[38;2;205;189;157mp[38;2;204;187;154mq[38;2;183;168;141mO[38;2;139;125;104mz[38;2;153;138;115mU[38;2;222;205;164mk[38;2;214;197;153md[38;2;207;196;168md[38;2;243;235;217mW[38;2;255;239;206mW[38;2;214;200;170mb[38;2;42;39;36ml[38;2;0;0;0m                            [38;2;0;0;0m");
  $display("[38;2;73;64;30m+[38;2;235;209;102mq[38;2;251;216;85mp[38;2;252;217;85mp[38;2;251;220;85mp[38;2;250;220;85mp[38;2;250;221;85mp[38;2;253;225;87md[38;2;254;229;91md[38;2;255;230;98mb[38;2;255;231;105mk[38;2;254;232;110mk[38;2;253;233;116mk[38;2;252;234;127mh[38;2;252;238;144mo[38;2;254;244;162m#[38;2;255;242;162m*[38;2;253;239;142mo[38;2;244;225;106md[38;2;245;218;87mp[38;2;245;215;95mp[38;2;174;142;64mX[38;2;204;178;88m0[38;2;235;211;93mq[38;2;216;188;95mZ[38;2;163;136;64mz[38;2;212;187;94mO[38;2;247;218;89mp[38;2;246;216;91mp[38;2;251;227;107mb[38;2;253;234;115mk[38;2;252;235;119mh[38;2;251;236;128mh[38;2;251;238;145mo[38;2;252;241;162m*[38;2;200;184;112mZ[38;2;197;176;81mQ[38;2;228;205;103mw[38;2;154;126;63mv[38;2;182;156;74mU[38;2;239;218;93mp[38;2;247;223;86mp[38;2;249;227;98md[38;2;253;232;115mk[38;2;253;233;122mh[38;2;254;235;121mh[38;2;253;235;117mk[38;2;247;228;100md[38;2;247;218;90mp[38;2;252;221;98md[38;2;188;166;89mL[38;2;37;29;18m;[38;2;0;0;2m [38;2;1;1;1m  [38;2;0;0;0m                           [38;2;1;1;1m  [38;2;0;0;0m [38;2;17;16;15m^[38;2;136;134;129mU[38;2;212;206;189mh[38;2;247;237;208mW[38;2;250;236;202mW[38;2;253;238;204mW[38;2;225;211;178mh[38;2;224;210;177mh[38;2;254;239;205mW[38;2;252;236;202mW[38;2;252;236;203mW[38;2;226;210;176mh[38;2;213;197;163md[38;2;249;236;198mM[38;2;253;239;202mW[38;2;249;235;196mM[38;2;217;203;162mb[38;2;199;184;145mw[38;2;187;169;132mO[38;2;172;151;114mC[38;2;136;109;76mu[38;2;126;94;62mr[38;2;136;101;62mx[38;2;142;104;57mn[38;2;152;112;62mu[38;2;150;116;70mv[38;2;168;147;112mC[38;2;182;175;156mm[38;2;229;227;219mM[38;2;252;250;241m@[38;2;251;250;238mB[38;2;252;249;237mB[38;2;254;247;231mB[38;2;254;246;232mB[38;2;254;247;236mB[38;2;254;238;213m&[38;2;222;190;137mp[38;2;231;187;119mq[38;2;232;185;114mw[38;2;230;182;114mw[38;2;229;181;112mw[38;2;227;181;112mm[38;2;232;184;118mw[38;2;238;189;121mq[38;2;244;198;131md[38;2;230;194;140md[38;2;80;57;36m+[38;2;113;99;87mx[38;2;189;181;157mw[38;2;178;166;143mO[38;2;199;184;154mq[38;2;173;158;128mQ[38;2;137;120;99mc[38;2;143;126;109mX[38;2;131;112;86mu[38;2;186;163;122m0[38;2;251;236;197mM[38;2;255;249;226mB[38;2;252;241;214m&[38;2;234;220;187mo[38;2;56;52;42mi[38;2;0;1;2m [38;2;0;0;0m                           [38;2;0;0;0m");
  $display("[38;2;72;66;29m+[38;2;232;210;101mq[38;2;250;216;84mp[38;2;251;217;84mp[38;2;250;220;84mp[38;2;249;220;84mp[38;2;249;219;84mp[38;2;250;221;84mp[38;2;250;224;86mp[38;2;251;226;89md[38;2;252;229;89md[38;2;250;229;95md[38;2;252;232;111mk[38;2;254;234;122mh[38;2;251;235;132ma[38;2;254;241;153m*[38;2;254;244;165m#[38;2;255;244;159m*[38;2;251;235;131mh[38;2;246;217;94mp[38;2;249;220;89mp[38;2;218;193;92mZ[38;2;149;127;61mv[38;2;229;200;99mw[38;2;235;205;93mw[38;2;207;187;97mO[38;2;127;103;54mr[38;2;225;196;92mm[38;2;248;218;87mp[38;2;242;218;91mp[38;2;246;228;105mb[38;2;251;233;119mk[38;2;253;234;122mh[38;2;252;236;129mh[38;2;252;239;139ma[38;2;254;243;148m*[38;2;206;188;95mO[38;2;217;191;88mZ[38;2;241;215;104mp[38;2;156;132;64mc[38;2;165;139;62mz[38;2;246;220;91mp[38;2;246;224;83mp[38;2;249;228;99mb[38;2;254;234;113mk[38;2;255;234;117mh[38;2;255;235;123mh[38;2;253;235;118mh[38;2;250;225;97md[38;2;252;215;85mp[38;2;255;222;99mb[38;2;187;168;96mL[38;2;32;29;15m,[38;2;0;1;1m [38;2;1;1;3m [38;2;0;0;0m                          [38;2;1;1;1m  [38;2;0;0;0m [38;2;13;13;13m'[38;2;144;142;136mJ[38;2;219;215;202mo[38;2;246;239;218m&[38;2;248;237;208mW[38;2;251;238;206mW[38;2;236;223;191m*[38;2;224;208;177mh[38;2;255;238;204mW[38;2;251;235;198mM[38;2;247;232;192m#[38;2;237;221;181mo[38;2;236;221;179mo[38;2;251;236;195mM[38;2;252;236;195mM[38;2;245;229;188m#[38;2;217;201;160mb[38;2;182;167;126m0[38;2;170;154;116mC[38;2;166;148;113mC[38;2;139;117;81mv[38;2;122;93;54mj[38;2;136;101;60mx[38;2;154;119;76mc[38;2;158;120;80mz[38;2;134;96;58mx[38;2;122;88;58mj[38;2;130;110;94mv[38;2;139;132;126mY[38;2;212;210;203ma[38;2;253;250;241m@[38;2;252;250;238mB[38;2;251;249;234mB[38;2;254;246;231mB[38;2;254;247;233mB[38;2;241;234;216mW[38;2;164;146;119mC[38;2;210;173;113mZ[38;2;246;194;118mp[38;2;250;193;117mp[38;2;242;191;116mp[38;2;229;182;113mw[38;2;221;177;110mZ[38;2;209;165;97m0[38;2;227;180;107mm[38;2;244;194;116mp[38;2;244;199;128md[38;2;147;117;80mv[38;2;152;135;109mY[38;2;249;241;209mW[38;2;239;231;214mM[38;2;211;204;194mh[38;2;162;153;140mQ[38;2;110;101;89mx[38;2;61;53;43m~[38;2;132;119;93mv[38;2;248;226;173m*[38;2;240;220;173mo[38;2;245;233;207mM[38;2;254;246;236mB[38;2;247;232;212mW[38;2;134;130;109mX[38;2;10;11;11m'[38;2;3;4;6m [38;2;1;1;1m [38;2;0;0;0m                         [38;2;0;0;0m");
  $display("");
  $display("\033[1;0m");
endtask

endmodule