`define CYCLE_TIME_clk1 47.1
`define CYCLE_TIME_clk2 10.1

`define SEED_NUMBER 38503729
`define PATTERN_NUMBER 10

module PATTERN(
	output reg clk1, clk2, rst_n, in_valid,
  output reg [17:0] in_row,
  output reg [11:0] in_kernel,
  input out_valid,
  input [7:0] out_data
);
//================================================================
// clock
//================================================================
real CYCLE_clk1 = `CYCLE_TIME_clk1;
always #(CYCLE_clk1/2.0) clk1 = ~clk1;
real CYCLE_clk2 = `CYCLE_TIME_clk2;
always #(CYCLE_clk2/2.0) clk2 = ~clk2;
//================================================================
// parameters & integer
//================================================================
integer SEED;
integer pat_count;
integer i, j, k;
integer exe_latency, total_latency;
integer rec_count;
//================================================================
// wire & registers 
//================================================================
reg [2:0] test_mtx[0:5][0:5];
reg [2:0] test_knl[0:5][0:3];

reg [7:0] golden[0:5][0:4][0:4];
reg [7:0] rec_out[0:5][0:4][0:4];
reg check;
//================================================================
// Main flow
//================================================================
initial begin
  reset_task;
  for(pat_count = 0; pat_count < `PATTERN_NUMBER; pat_count = pat_count + 1) begin
    input_task;
    ans_gen_task;
    wait_task;
    check_task;
  end
  YOU_PASS_task;
end

always @(negedge clk1) begin
  if(out_valid === 1'b0 && out_data !== 8'd0) begin : OUT_RESET_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("      Output must be 0 when out_valid is low      ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk1);
    $finish;
  end
  if(in_valid === 1'b1 && out_valid === 1'b1) begin : OVERLAP_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("   in_valid and out_valid cannot be high at once  ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk1);
    $finish;
  end
end
//================================================================
// task
//================================================================
task reset_task;
  SEED = `SEED_NUMBER;
  rst_n = 1'b1;
  in_valid = 1'b0;
  in_row = 'dx; in_kernel = 'dx;

  total_latency = 0;

  force clk1 = 'b0; force clk2 = 'b0;
  #(CYCLE_clk1 * ($random(SEED) % 'd3 + 'd1)); rst_n = 'b0;
  #(CYCLE_clk1 * 0.75);

  if(out_valid !== 1'b0 || out_data !== 8'b0) begin : RESET_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("           Output must be 0 after reset           ");
    $display("--------------------------------------------------");
      #(CYCLE_clk1 * 5);
    $finish;
  end

  #(CYCLE_clk1 * 0.25); rst_n = 'b1;
  #(CYCLE_clk1); release clk1; release clk2;
  repeat(3) @(negedge clk1);
endtask

task input_task;
  repeat($random(SEED) % 'd3) @(negedge clk1);
  // Generate random inputs
  foreach(test_mtx[i, j]) test_mtx[i][j] = $random(SEED) % 'd8;
  foreach(test_knl[i, j]) test_knl[i][j] = $random(SEED) % 'd4;
  // Send inputs
  in_valid = 1'b1;
  for(i = 0; i < 6; i = i + 1) begin
    in_row = {test_mtx[i][5], test_mtx[i][4], test_mtx[i][3],
              test_mtx[i][2], test_mtx[i][1], test_mtx[i][0]};
    in_kernel = {test_knl[i][3], test_knl[i][2], test_knl[i][1], test_knl[i][0]};
      @(negedge clk1);
  end
  // Reset inputs
  in_valid = 1'b0;
  in_row = 'dx; in_kernel = 'dx;
    @(negedge clk1);
  exe_latency = 1;
endtask

task ans_gen_task;
  for(i = 0; i < 6; i = i + 1) begin
    for(j = 0; j < 5; j = j + 1) begin
      for(k = 0; k < 5; k = k + 1) begin
        golden[i][j][k] = 8'd0;
        golden[i][j][k] = golden[i][j][k] +     test_mtx[j][k] * test_knl[i][0];
        golden[i][j][k] = golden[i][j][k] +   test_mtx[j][k+1] * test_knl[i][1];
        golden[i][j][k] = golden[i][j][k] +   test_mtx[j+1][k] * test_knl[i][2];
        golden[i][j][k] = golden[i][j][k] + test_mtx[j+1][k+1] * test_knl[i][3];
      end
    end
  end
endtask

task wait_task;
  while(out_valid !== 1'b1) begin
    exe_latency = exe_latency + 1;
    if(exe_latency == 5000) begin : TIMEOUT_CHECK
      fail_task;
      $display("--------------------------------------------------");
      $display("                      FAIL!!                      ");
      $display("       Execution timeout (over 5000 cycles)       ");
      $display("--------------------------------------------------");
      repeat(5) @(negedge clk1);
      $finish;
    end
      @(negedge clk1);
  end
endtask

task check_task;
  i = 0; j = 0; k = 0;
  rec_count = 0;
  check = 1'b0;
  while(rec_count < 150) begin
    rec_count = rec_count + 1;
    rec_out[i][j][k] = out_data;
    check = check || (rec_out[i][j][k] !== golden[i][j][k]);
      @(negedge clk1);
    exe_latency = exe_latency + 1;
    if(rec_count != 150)
      wait_task;
    k = (k + 1) % 5;
    j = (j + (k == 0)) % 5;
    i = (i + (j == 0 && k == 0)) % 6;
  end
    @(negedge clk1);
  if(out_valid !== 1'b0) begin
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("        out_valid must be low after output        ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk1);
    $finish;
  end
  if(check) begin
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("         Output does not match with golden        ");
    $display("==================================================");
    $display("  Input Matrix:");
    for(i = 0; i < 6; i = i + 1) begin
      $write("                ");
      for(j = 0; j < 6; j = j + 1) begin
        $write(" %1d", test_mtx[i][j]);
      end
      $display("");
    end
    $display("  Kernel Matrix:");
    for(i = 0; i < 2; i = i + 1) begin
      $write("     ");
      for(j = 0; j < 6; j = j + 1) begin
        $write(" %1d %1d |", test_knl[j][i*2], test_knl[j][i*2+1]);
      end
      $display("");
    end
    $display("--------------------------------------------------");
    $display("  Golden:");
    for(i = 0; i < 5; i = i + 1) begin
      for(j = 0; j < 6; j = j + 1) begin
        for(k = 0; k < 5; k = k + 1) begin
          $write(" %3d", golden[j][i][k]);
        end
        $write(" |");
      end
      $display("");
    end
    $display("\n  Yours:");
    for(i = 0; i < 5; i = i + 1) begin
      for(j = 0; j < 6; j = j + 1) begin
        for(k = 0; k < 5; k = k + 1) begin
          if(rec_out[j][i][k] !== golden[j][i][k])
            $write("\033[38;5;196m %3d\033[0m", rec_out[j][i][k]);
          else
            $write(" %3d", rec_out[j][i][k]);
        end
        $write(" |");
      end
      $display("");
    end
    $display("\n--------------------------------------------------");
    repeat(5) @(negedge clk1);
    $finish;
  end
  $display("\033[38;5;123mPATTERN NO.%4d PASS!!\033[0;32m EXECUTION CYCLE :%4d\033[m", pat_count, exe_latency);
  total_latency = total_latency + exe_latency;
endtask

task YOU_PASS_task;
  $display("\033[38;2;255;255;255m                                                                                    \033[38;2;255;255;254m \033[38;2;255;255;255m                                   ");
  $display("\033[38;2;255;255;255m                                                                                  \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;246;243;240mB\033[38;2;226;223;208m#\033[38;2;231;232;224mW\033[38;2;236;237;233m&\033[38;2;255;255;255m                                ");
  $display("\033[38;2;255;255;255m                                                                                    \033[38;2;254;254;252m \033[38;2;228;227;215mM\033[38;2;209;211;190mh\033[38;2;188;197;178md\033[38;2;172;177;169mw\033[38;2;210;208;207ma\033[38;2;254;253;251m \033[38;2;255;255;255m  \033[38;2;255;255;254m \033[38;2;255;255;255m                          ");
  $display("\033[38;2;255;255;255m                                                                                     \033[38;2;254;254;252m \033[38;2;223;222;209m*\033[38;2;235;236;215mW\033[38;2;224;235;212mM\033[38;2;148;168;152m0\033[38;2;114;130;126mX\033[38;2;194;199;199mk\033[38;2;255;255;255m                            ");
  $display("\033[38;2;255;255;255m                                                           \033[38;2;254;255;255m  \033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;255;255;255m          \033[38;2;254;255;255m \033[38;2;255;255;255m            \033[38;2;246;245;243mB\033[38;2;198;198;179mb\033[38;2;239;249;223m&\033[38;2;173;196;177mp\033[38;2;136;170;155m0\033[38;2;85;118;106mu\033[38;2;117;133;127mY\033[38;2;229;229;227mW\033[38;2;255;255;255m   \033[38;2;254;255;255m \033[38;2;255;255;255m   \033[38;2;254;255;255m  \033[38;2;255;255;255m                 ");
  $display("\033[38;2;255;255;255m                                                          \033[38;2;254;255;255m \033[38;2;254;253;255m \033[38;2;249;253;252m@\033[38;2;250;254;254m \033[38;2;255;255;255m      \033[38;2;254;254;251m \033[38;2;244;244;240mB\033[38;2;246;247;244mB\033[38;2;253;252;252m \033[38;2;255;255;255m               \033[38;2;212;212;201ma\033[38;2;212;216;195ma\033[38;2;204;212;191mh\033[38;2;237;245;220m&\033[38;2;213;236;215m#\033[38;2;138;164;149mQ\033[38;2;86;98;90mx\033[38;2;194;193;193mb\033[38;2;255;255;255m \033[38;2;254;255;255m  \033[38;2;255;255;255m   \033[38;2;253;255;254m \033[38;2;254;255;254m \033[38;2;230;233;229mW\033[38;2;205;214;208mo\033[38;2;254;254;253m \033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                                                          \033[38;2;254;255;254m \033[38;2;255;254;254m \033[38;2;220;244;237m&\033[38;2;152;230;211mk\033[38;2;198;237;228m#\033[38;2;232;245;235m&\033[38;2;248;252;248m@\033[38;2;254;255;255m \033[38;2;255;255;255m  \033[38;2;253;253;252m \033[38;2;210;211;206mo\033[38;2;124;133;126mY\033[38;2;84;108;101mn\033[38;2;101;132;126mX\033[38;2;116;140;136mU\033[38;2;129;147;143mC\033[38;2;137;153;149mL\033[38;2;147;159;157m0\033[38;2;162;170;169mm\033[38;2;176;178;177mq\033[38;2;189;189;189md\033[38;2;211;211;210mo\033[38;2;247;246;245mB\033[38;2;255;255;255m   \033[38;2;255;254;255m \033[38;2;255;255;255m \033[38;2;245;243;239mB\033[38;2;182;182;167mq\033[38;2;224;231;206m#\033[38;2;239;248;226m&\033[38;2;141;168;151m0\033[38;2;100;147;129mY\033[38;2;130;164;151mQ\033[38;2;81;97;92mr\033[38;2;192;191;189mb\033[38;2;255;255;255m \033[38;2;255;253;255m \033[38;2;255;255;255m   \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;217;224;218m#\033[38;2;93;124;113mc\033[38;2;123;151;143mC\033[38;2;220;222;221m#\033[38;2;255;255;255m \033[38;2;253;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                           \033[38;2;255;254;254m \033[38;2;248;254;253m@\033[38;2;165;231;218ma\033[38;2;139;222;200md\033[38;2;215;237;224mM\033[38;2;210;232;220m#\033[38;2;204;232;218m*\033[38;2;229;240;233m&\033[38;2;243;249;246mB\033[38;2;253;255;253m \033[38;2;255;255;255m \033[38;2;239;240;239m8\033[38;2;136;148;145mL\033[38;2;36;73;65m_\033[38;2;32;90;78m-\033[38;2;30;92;81m?\033[38;2;29;88;79m-\033[38;2;30;85;78m-\033[38;2;32;82;77m-\033[38;2;30;78;72m_\033[38;2;30;70;65m+\033[38;2;31;60;54m~\033[38;2;62;82;76m1\033[38;2;144;156;149mQ\033[38;2;219;226;221m#\033[38;2;254;255;255m \033[38;2;255;255;255m  \033[38;2;255;255;254m \033[38;2;174;173;162mm\033[38;2;228;235;211mM\033[38;2;226;234;213mM\033[38;2;198;212;193mh\033[38;2;138;178;163mO\033[38;2;48;111;101mr\033[38;2;68;115;111mn\033[38;2;96;115;111mv\033[38;2;240;240;239m8\033[38;2;255;254;255m \033[38;2;255;255;255m     \033[38;2;242;245;241mB\033[38;2;141;163;149mQ\033[38;2;149;188;170mm\033[38;2;82;110;101mn\033[38;2;198;202;201mh\033[38;2;255;255;255m \033[38;2;253;255;255m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                           \033[38;2;254;254;254m \033[38;2;254;255;255m \033[38;2;246;251;251m@\033[38;2;163;231;215mh\033[38;2;179;237;227m*\033[38;2;253;255;253m \033[38;2;252;255;250m \033[38;2;239;251;244mB\033[38;2;221;243;233mW\033[38;2;220;242;231mW\033[38;2;231;248;239m8\033[38;2;251;255;255m \033[38;2;255;255;255m \033[38;2;174;177;173mw\033[38;2;51;77;73m?\033[38;2;43;95;89m1\033[38;2;39;97;89m1\033[38;2;41;96;88m1\033[38;2;39;95;86m1\033[38;2;37;96;87m1\033[38;2;38;96;89m1\033[38;2;37;95;88m1\033[38;2;29;87;77m-\033[38;2;19;72;62m~\033[38;2;42;91;82m?\033[38;2;99;137;129mX\033[38;2;164;190;184mq\033[38;2;214;225;223m#\033[38;2;249;250;251m@\033[38;2;172;170;161mm\033[38;2;204;210;189mh\033[38;2;206;213;193ma\033[38;2;233;243;215mW\033[38;2;240;251;227m8\033[38;2;157;192;179mq\033[38;2;41;101;97mf\033[38;2;48;90;86m1\033[38;2;200;203;200mh\033[38;2;255;255;255m      \033[38;2;241;243;240m8\033[38;2;158;166;149mO\033[38;2;225;242;222mW\033[38;2;110;147;130mU\033[38;2;60;96;86mf\033[38;2;218;217;219m*\033[38;2;255;255;255m           ");
  $display("\033[38;2;255;255;255m                                                              \033[38;2;240;241;241m8\033[38;2;149;213;203md\033[38;2;154;228;221mh\033[38;2;166;182;182mq\033[38;2;148;147;145mL\033[38;2;150;150;148mQ\033[38;2;162;163;158mO\033[38;2;169;183;171mw\033[38;2;176;200;189md\033[38;2;209;226;221m*\033[38;2;252;255;255m \033[38;2;151;159;155m0\033[38;2;38;73;65m_\033[38;2;40;97;84m1\033[38;2;41;96;85m1\033[38;2;39;97;87m1\033[38;2;38;97;89m1\033[38;2;38;95;88m1\033[38;2;38;95;86m1\033[38;2;37;96;84m1\033[38;2;33;98;84m?\033[38;2;28;86;75m-\033[38;2;17;64;56mi\033[38;2;20;62;56mi\033[38;2;44;108;105mj\033[38;2;99;166;162mC\033[38;2;90;106;103mn\033[38;2;191;197;179md\033[38;2;234;243;221mW\033[38;2;235;244;221m&\033[38;2;237;246;222m&\033[38;2;237;249;227m&\033[38;2;143;186;171mm\033[38;2;32;80;73m_\033[38;2;129;138;133mJ\033[38;2;255;255;255m      \033[38;2;224;226;223mM\033[38;2;156;162;148m0\033[38;2;207;214;191ma\033[38;2;186;209;183mb\033[38;2;93;159;144mU\033[38;2;98;138;136mY\033[38;2;247;247;247m@\033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                         \033[38;2;245;244;244mB\033[38;2;219;219;218m*\033[38;2;183;187;184mp\033[38;2;139;150;147mL\033[38;2;94;114;110mv\033[38;2;65;92;87mj\033[38;2;48;88;81m1\033[38;2;41;163;152mz\033[38;2;45;173;171mU\033[38;2;23;102;97m1\033[38;2;20;70;63m~\033[38;2;25;60;53mi\033[38;2;27;47;41m!\033[38;2;23;30;26m;\033[38;2;25;27;29m;\033[38;2;56;77;79m?\033[38;2;87;126;123mc\033[38;2;38;92;89m1\033[38;2;43;130;121mn\033[38;2;37;121;114mr\033[38;2;39;104;99mf\033[38;2;39;97;92mf\033[38;2;40;97;88m1\033[38;2;38;96;84m1\033[38;2;38;95;86m1\033[38;2;38;95;85m1\033[38;2;35;96;84m?\033[38;2;37;93;83m?\033[38;2;23;63;58m~\033[38;2;3;23;20m \033[38;2;10;32;33m;\033[38;2;44;64;60m+\033[38;2;223;231;213m#\033[38;2;237;248;224m&\033[38;2;235;243;223m&\033[38;2;237;243;223m&\033[38;2;240;245;220m&\033[38;2;219;239;217mM\033[38;2;97;146;133mY\033[38;2;81;102;95mx\033[38;2;250;248;247m@\033[38;2;255;255;255m   \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;180;180;175mq\033[38;2;161;164;148mO\033[38;2;217;224;201m*\033[38;2;202;216;196ma\033[38;2;110;169;152mL\033[38;2;50;157;143mz\033[38;2;177;199;197mb\033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                     \033[38;2;246;247;247mB\033[38;2;208;213;210mo\033[38;2;162;173;169mm\033[38;2;108;126;123mX\033[38;2;71;99;96mr\033[38;2;49;89;83m1\033[38;2;39;90;80m?\033[38;2;37;94;84m?\033[38;2;35;99;89m1\033[38;2;35;105;91mf\033[38;2;45;102;91mf\033[38;2;39;104;97mf\033[38;2;40;156;145mc\033[38;2;55;201;191mQ\033[38;2;51;180;174mJ\033[38;2;40;144;135mv\033[38;2;38;114;101mj\033[38;2;44;90;82m1\033[38;2;15;34;35m;\033[38;2;0;0;0m \033[38;2;1;3;4m \033[38;2;12;29;29m,\033[38;2;39;108;102mj\033[38;2;44;143;134mv\033[38;2;49;139;131mv\033[38;2;40;103;95mf\033[38;2;41;97;88m1\033[38;2;40;97;88m1\033[38;2;38;95;86m1\033[38;2;39;95;87m1\033[38;2;38;95;86m1\033[38;2;37;95;86m1\033[38;2;37;94;84m?\033[38;2;23;54;50m!\033[38;2;0;0;0m \033[38;2;120;123;115mX\033[38;2;245;251;233mB\033[38;2;235;245;221m&\033[38;2;240;243;222m&\033[38;2;242;243;222m&\033[38;2;236;244;221m&\033[38;2;238;244;223m&\033[38;2;165;198;181mp\033[38;2;67;89;81mf\033[38;2;232;228;227mW\033[38;2;255;255;255m    \033[38;2;244;244;242mB\033[38;2;131;132;123mU\033[38;2;211;215;198ma\033[38;2;212;219;196mo\033[38;2;199;212;191mh\033[38;2;186;230;205ma\033[38;2;55;189;176mC\033[38;2;124;172;169m0\033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m       ");
  $display("\033[38;2;255;255;255m                                                   \033[38;2;238;240;237m8\033[38;2;160;165;159mO\033[38;2;89;106;99mn\033[38;2;47;79;72m-\033[38;2;36;82;73m-\033[38;2;32;90;79m?\033[38;2;37;102;91mf\033[38;2;44;110;98mj\033[38;2;47;111;98mj\033[38;2;48;110;99mj\033[38;2;46;108;97mj\033[38;2;45;107;95mj\033[38;2;42;110;96mj\033[38;2;40;117;108mr\033[38;2;27;146;136mu\033[38;2;50;203;192mQ\033[38;2;100;251;247mk\033[38;2;54;202;193mQ\033[38;2;30;131;121mx\033[38;2;40;106;95mf\033[38;2;44;91;83m1\033[38;2;10;25;24m,\033[38;2;1;0;1m \033[38;2;2;0;1m \033[38;2;32;60;55m~\033[38;2;45;100;88mf\033[38;2;41;98;90mf\033[38;2;40;100;91mf\033[38;2;41;99;90mf\033[38;2;41;98;90mf\033[38;2;40;97;88m1\033[38;2;41;97;88m1\033[38;2;38;95;86m1\033[38;2;37;95;86m1\033[38;2;40;97;87m1\033[38;2;21;58;50mi\033[38;2;56;63;54m_\033[38;2;221;226;207m*\033[38;2;239;249;227m8\033[38;2;236;246;222m&\033[38;2;232;237;215mW\033[38;2;221;225;203m*\033[38;2;236;244;221m&\033[38;2;239;242;222m&\033[38;2;210;231;210m*\033[38;2;88;114;100mu\033[38;2;93;110;106mu\033[38;2;171;183;182mq\033[38;2;243;243;243mB\033[38;2;255;255;255m  \033[38;2;166;164;159mZ\033[38;2;167;170;156mZ\033[38;2;218;223;203m*\033[38;2;223;228;203m*\033[38;2;231;246;223m&\033[38;2;148;212;194mp\033[38;2;44;194;190mC\033[38;2;127;178;178mO\033[38;2;255;255;255m  \033[38;2;255;254;255m \033[38;2;255;255;255m       ");
  $display("\033[38;2;255;255;255m                                                   \033[38;2;247;247;244mB\033[38;2;226;227;224mM\033[38;2;219;220;217m*\033[38;2;202;205;202mh\033[38;2;175;182;180mq\033[38;2;134;148;145mC\033[38;2;87;108;105mu\033[38;2;51;83;78m?\033[38;2;34;84;74m-\033[38;2;41;102;90mf\033[38;2;47;111;99mj\033[38;2;45;110;100mj\033[38;2;34;131;119mx\033[38;2;52;192;181mC\033[38;2;78;235;233mp\033[38;2;90;236;236md\033[38;2;72;217;210mm\033[38;2;34;157;149mc\033[38;2;37;115;102mj\033[38;2;41;105;91mf\033[38;2;43;107;94mj\033[38;2;22;53;47m!\033[38;2;1;1;3m \033[38;2;1;0;1m \033[38;2;25;51;46m!\033[38;2;47;105;94mj\033[38;2;42;102;92mf\033[38;2;43;100;91mff\033[38;2;44;100;91mf\033[38;2;43;98;90mf\033[38;2;41;97;90mf\033[38;2;38;91;84m?\033[38;2;33;77;71m_\033[38;2;35;67;63m+\033[38;2;90;105;96mn\033[38;2;220;225;209m*\033[38;2;245;250;227m8\033[38;2;237;248;224m&\033[38;2;234;244;220mW\033[38;2;206;213;190mh\033[38;2;216;224;201mo\033[38;2;222;232;208m#\033[38;2;237;243;220m&\033[38;2;233;244;222m&\033[38;2;142;168;151m0\033[38;2;16;45;41ml\033[38;2;41;106;100mj\033[38;2;108;141;137mU\033[38;2;229;229;229mW\033[38;2;188;185;181mp\033[38;2;154;154;143mQ\033[38;2;232;240;218mW\033[38;2;231;240;217mW\033[38;2;233;240;218mW\033[38;2;205;238;215m#\033[38;2;73;202;190m0\033[38;2;49;184;177mJ\033[38;2;193;206;206mh\033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                          \033[38;2;225;221;222m#\033[38;2;155;154;155m0\033[38;2;74;87;84mj\033[38;2;34;65;57m~\033[38;2;41;91;81m?\033[38;2;41;132;120mn\033[38;2;46;175;165mU\033[38;2;50;181;173mJ\033[38;2;41;153;144mc\033[38;2;34;131;120mn\033[38;2;42;113;105mr\033[38;2;47;107;96mj\033[38;2;43;108;95mj\033[38;2;42;110;96mj\033[38;2;35;76;66m_\033[38;2;2;5;5m \033[38;2;1;0;0m \033[38;2;28;55;52mi\033[38;2;46;104;98mj\033[38;2;43;102;91mf\033[38;2;45;101;89mf\033[38;2;42;94;83m1\033[38;2;42;85;77m?\033[38;2;37;77;69m_\033[38;2;44;76;69m-\033[38;2;71;91;84mj\033[38;2;120;129;120mX\033[38;2;188;194;181md\033[38;2;239;246;226m&\033[38;2;243;250;225m8\033[38;2;239;246;222m&\033[38;2;226;234;212mM\033[38;2;213;221;198mo\033[38;2;236;237;216mW\033[38;2;242;244;223m&\033[38;2;225;235;211mM\033[38;2;214;220;198mo\033[38;2;241;246;224m&\033[38;2;203;218;200ma\033[38;2;44;52;44mi\033[38;2;1;18;16m'\033[38;2;47;125;119mn\033[38;2;66;102;101mr\033[38;2;139;147;134mC\033[38;2;232;240;218mW\033[38;2;234;241;217mW\033[38;2;232;240;218mW\033[38;2;226;243;220mW\033[38;2;128;210;195mq\033[38;2;45;188;183mC\033[38;2;138;185;184mm\033[38;2;255;253;252m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                  \033[38;2;254;255;255m \033[38;2;255;255;255m   \033[38;2;252;251;251m@\033[38;2;226;228;227mM\033[38;2;187;199;196mb\033[38;2;158;171;168mZ\033[38;2;155;165;162mO\033[38;2;155;167;162mO\033[38;2;132;142;139mJ\033[38;2;44;55;53m~\033[38;2;25;46;41ml\033[38;2;32;71;64m+\033[38;2;36;92;85m?\033[38;2;46;110;99mj\033[38;2;42;101;88mf\033[38;2;48;104;91mj\033[38;2;50;109;98mj\033[38;2;48;110;99mj\033[38;2;46;109;100mj\033[38;2;45;110;98mj\033[38;2;48;101;90mf\033[38;2;21;44;39ml\033[38;2;0;1;2m \033[38;2;31;55;53mi\033[38;2;50;105;99mj\033[38;2;42;102;93mf\033[38;2;44;104;91mf\033[38;2;42;89;79m?\033[38;2;61;73;69m?\033[38;2;178;183;171mq\033[38;2;211;218;200mo\033[38;2;235;242;221mW\033[38;2;249;255;233mB\033[38;2;246;254;230mB\033[38;2;237;246;222m&\033[38;2;230;239;215mW\033[38;2;215;223;200mo\033[38;2;216;224;201mo\033[38;2;234;243;220mW\033[38;2;241;243;222m&\033[38;2;240;243;222m&\033[38;2;237;244;222m&\033[38;2;213;223;200mo\033[38;2;228;235;209mM\033[38;2;235;248;226m&\033[38;2;114;129;116mX\033[38;2;0;0;0m \033[38;2;20;32;34m;\033[38;2;133;151;143mC\033[38;2;231;243;225m&\033[38;2;236;241;220mW\033[38;2;233;239;215mW\033[38;2;231;245;221mW\033[38;2;181;233;214mo\033[38;2;56;183;170mJ\033[38;2;101;160;157mC\033[38;2;244;241;239m8\033[38;2;254;255;255m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                   \033[38;2;244;244;241mB\033[38;2;203;209;206ma\033[38;2;145;164;160m0\033[38;2;97;130;122mz\033[38;2;64;110;99mx\033[38;2;45;103;90mf\033[38;2;41;100;87mf\033[38;2;43;99;88mf\033[38;2;42;99;88mf\033[38;2;42;103;92mf\033[38;2;53;118;108mx\033[38;2;51;114;104mr\033[38;2;52;103;92mj\033[38;2;43;71;64m_\033[38;2;28;50;45m!\033[38;2;42;76;69m-\033[38;2;45;91;82m1\033[38;2;49;109;98mj\033[38;2;47;108;98mj\033[38;2;48;106;98mj\033[38;2;46;107;96mj\033[38;2;47;108;97mj\033[38;2;51;103;96mj\033[38;2;33;66;63m+\033[38;2;9;27;24m,\033[38;2;34;65;59m~\033[38;2;41;96;85m1\033[38;2;35;92;80m?\033[38;2;38;84;76m-\033[38;2;33;49;43m!\033[38;2;107;112;99mv\033[38;2;216;222;202mo\033[38;2;241;249;227m8\033[38;2;238;246;223m&\033[38;2;227;235;211mM\033[38;2;222;230;207m#\033[38;2;228;236;213mM\033[38;2;235;242;220mW\033[38;2;240;248;224m&\033[38;2;238;247;223m&\033[38;2;240;243;222m&\033[38;2;241;243;222m&\033[38;2;238;244;222m&\033[38;2;223;236;211mM\033[38;2;193;205;180mb\033[38;2;238;251;226m8\033[38;2;196;209;189mk\033[38;2;24;42;34mI\033[38;2;105;128;119mz\033[38;2;231;243;226m&\033[38;2;224;224;203m*\033[38;2;228;234;211mM\033[38;2;234;244;220mW\033[38;2;199;244;226mM\033[38;2;89;204;187mO\033[38;2;80;151;147mY\033[38;2;230;232;230mW\033[38;2;255;255;254m \033[38;2;253;255;254m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                                \033[38;2;248;249;249m@\033[38;2;203;212;210ma\033[38;2;142;163;157m0\033[38;2;85;121;112mv\033[38;2;53;105;93mj\033[38;2;43;105;94mf\033[38;2;46;110;99mj\033[38;2;50;112;100mr\033[38;2;47;115;104mr\033[38;2;54;150;131mc\033[38;2;51;141;124mv\033[38;2;48;112;100mr\033[38;2;49;115;103mr\033[38;2;50;118;105mx\033[38;2;46;114;103mr\033[38;2;52;112;102mr\033[38;2;57;114;101mr\033[38;2;36;68;61m+\033[38;2;7;12;13m'\033[38;2;22;40;38mI\033[38;2;47;99;89mf\033[38;2;47;108;99mj\033[38;2;48;105;97mj\033[38;2;46;106;96mjj\033[38;2;46;105;96mj\033[38;2;47;107;96mj\033[38;2;43;90;79m?\033[38;2;29;47;41m!\033[38;2;76;92;85mj\033[38;2;126;143;130mJ\033[38;2;161;173;156mZ\033[38;2;190;197;181md\033[38;2;185;192;179md\033[38;2;125;136;123mU\033[38;2;138;149;134mC\033[38;2;211;221;204mo\033[38;2;243;252;233mB\033[38;2;247;255;234mB\033[38;2;242;252;228m8\033[38;2;239;249;224m&\033[38;2;240;249;224m&\033[38;2;239;248;225m&\033[38;2;239;246;224m&\033[38;2;238;246;223m&\033[38;2;238;246;222m&\033[38;2;235;247;224m&\033[38;2;176;194;173mp\033[38;2;217;230;209m*\033[38;2;241;250;228m8\033[38;2;130;146;129mJ\033[38;2;81;96;86mr\033[38;2;196;203;188mk\033[38;2;219;222;201m*\033[38;2;239;244;222m&\033[38;2;190;232;212mo\033[38;2;91;203;189mO\033[38;2;58;130;125mu\033[38;2;212;216;214m*\033[38;2;255;255;255m \033[38;2;254;254;255m \033[38;2;254;255;254m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                              \033[38;2;242;242;241m8\033[38;2;177;185;176mq\033[38;2;102;126;115mz\033[38;2;52;95;82mf\033[38;2;39;93;79m?\033[38;2;40;100;90mf\033[38;2;46;111;100mj\033[38;2;51;116;105mr\033[38;2;51;116;104mr\033[38;2;51;113;100mr\033[38;2;46;110;98mj\033[38;2;48;125;109mx\033[38;2;51;120;107mx\033[38;2;52;113;103mr\033[38;2;52;114;103mr\033[38;2;52;113;102mr\033[38;2;50;113;102mr\033[38;2;52;112;102mr\033[38;2;51;113;102mr\033[38;2;55;111;102mr\033[38;2;21;42;38mI\033[38;2;0;0;0m \033[38;2;31;57;52mi\033[38;2;56;113;101mr\033[38;2;49;109;99mjj\033[38;2;48;108;98mjj\033[38;2;46;100;92mf\033[38;2;45;90;80m?\033[38;2;132;146;137mC\033[38;2;223;223;210m*\033[38;2;255;255;244m@\033[38;2;253;255;234m@\033[38;2;246;255;229mB\033[38;2;235;253;229m8\033[38;2;210;236;217m#\033[38;2;130;171;155m0\033[38;2;73;115;101mn\033[38;2;108;134;120mX\033[38;2;194;211;196mh\033[38;2;235;250;232m8\033[38;2;242;255;232mB\033[38;2;237;252;226m8\033[38;2;236;253;227m8\033[38;2;238;252;227m8\033[38;2;237;248;224m&\033[38;2;237;247;223m&\033[38;2;237;250;227m8\033[38;2;170;189;169mq\033[38;2;185;200;179md\033[38;2;234;240;218mW\033[38;2;234;237;217mW\033[38;2;208;211;193ma\033[38;2;231;237;219mW\033[38;2;228;238;217mM\033[38;2;149;192;170mm\033[38;2;56;158;148mX\033[38;2;40;145;139mv\033[38;2;154;163;165mO\033[38;2;255;255;255m  \033[38;2;254;255;255m  \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                                              \033[38;2;247;248;247m@\033[38;2;229;230;228mW\033[38;2;223;227;224mM\033[38;2;212;216;212mo\033[38;2;177;183;177mq\033[38;2;131;143;136mJ\033[38;2;85;103;96mx\033[38;2;51;82;75m?\033[38;2;41;85;77m?\033[38;2;51;103;93mj\033[38;2;52;113;100mr\033[38;2;45;110;96mj\033[38;2;51;114;99mr\033[38;2;51;114;101mr\033[38;2;53;112;105mr\033[38;2;52;113;105mr\033[38;2;51;115;103mr\033[38;2;51;113;102mr\033[38;2;49;114;102mr\033[38;2;54;117;106mx\033[38;2;45;84;78m?\033[38;2;1;5;6m \033[38;2;12;18;19m \033[38;2;57;101;93mj\033[38;2;50;114;102mr\033[38;2;50;111;100mr\033[38;2;50;109;100mr\033[38;2;47;105;97mj\033[38;2;41;93;87m1\033[38;2;44;94;86m1\033[38;2;48;104;91mj\033[38;2;57;98;87mf\033[38;2;136;153;138mC\033[38;2;233;242;221mW\033[38;2;245;252;229mB\033[38;2;237;247;226m&\033[38;2;221;241;223mW\033[38;2;149;204;186mq\033[38;2;62;134;114mu\033[38;2;27;65;49mi\033[38;2;11;31;18m,\033[38;2;78;107;90mx\033[38;2;198;229;209mo\033[38;2;244;255;235mB\033[38;2;240;252;229m8\033[38;2;239;251;227m8\033[38;2;238;248;225m&\033[38;2;238;246;223m&\033[38;2;238;250;226m8\033[38;2;186;206;185mb\033[38;2;170;183;162mw\033[38;2;238;239;218mW\033[38;2;239;242;220m&\033[38;2;226;235;213mM\033[38;2;201;218;198ma\033[38;2;153;176;158mZ\033[38;2;114;171;153mL\033[38;2;56;200;188mQ\033[38;2;46;123;124mn\033[38;2;224;218;213m*\033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                                               \033[38;2;245;243;244mB\033[38;2;215;216;216m*\033[38;2;182;188;186md\033[38;2;157;167;165mZ\033[38;2;136;150;145mL\033[38;2;120;133;129mY\033[38;2;76;86;84mj\033[38;2;15;22;23m,\033[38;2;9;16;18m'\033[38;2;23;38;37mI\033[38;2;30;63;57m~\033[38;2;45;99;85mf\033[38;2;53;119;105mx\033[38;2;49;114;106mr\033[38;2;50;115;106mr\033[38;2;47;109;97mj\033[38;2;48;112;97mj\033[38;2;49;116;100mr\033[38;2;50;116;100mr\033[38;2;53;102;90mj\033[38;2;6;18;14m'\033[38;2;1;3;3m \033[38;2;42;79;72m-\033[38;2;54;113;105mr\033[38;2;48;110;102mr\033[38;2;47;111;100mr\033[38;2;48;105;94mj\033[38;2;30;68;64m+\033[38;2;32;78;70m_\033[38;2;61;109;96mr\033[38;2;104;137;126mX\033[38;2;57;80;71m?\033[38;2;74;88;78mf\033[38;2;227;233;218mM\033[38;2;244;252;228m8\033[38;2;235;251;228m8\033[38;2;174;223;206mh\033[38;2;84;169;144mU\033[38;2;31;101;66m-\033[38;2;3;59;25mI\033[38;2;46;149;117mu\033[38;2;77;184;153mC\033[38;2;194;233;212mo\033[38;2;247;255;240m@\033[38;2;241;251;233m8\033[38;2;237;249;225m&\033[38;2;236;247;221m&\033[38;2;236;248;227m&\033[38;2;152;179;163mZ\033[38;2;147;164;148m0\033[38;2;245;245;226m8\033[38;2;225;232;209m#\033[38;2;187;197;176md\033[38;2;178;190;170mq\033[38;2;222;233;211m#\033[38;2;203;238;215m*\033[38;2;72;207;193mO\033[38;2;37;133;131mu\033[38;2;196;193;190mb\033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                                           \033[38;2;246;245;245mB\033[38;2;212;215;214mo\033[38;2;162;173;169mm\033[38;2;118;135;129mY\033[38;2;82;108;100mn\033[38;2;57;97;86mf\033[38;2;50;104;89mj\033[38;2;51;108;95mj\033[38;2;50;109;99mr\033[38;2;51;112;99mr\033[38;2;56;116;102mx\033[38;2;57;112;98mr\033[38;2;46;91;80m1\033[38;2;25;49;44m!\033[38;2;3;3;6m \033[38;2;26;46;42m!\033[38;2;60;118;104mx\033[38;2;52;118;106mx\033[38;2;55;116;105mx\033[38;2;44;96;85m1\033[38;2;22;61;52mi\033[38;2;52;106;92mj\033[38;2;56;115;99mr\033[38;2;33;63;56m~\033[38;2;2;5;4m \033[38;2;2;0;0m \033[38;2;28;54;51mi\033[38;2;57;113;105mx\033[38;2;49;111;103mr\033[38;2;47;111;101mr\033[38;2;51;109;96mj\033[38;2;41;75;63m_\033[38;2;74;103;87mr\033[38;2;186;201;184mb\033[38;2;242;246;232m8\033[38;2;165;179;163mm\033[38;2;119;128;120mX\033[38;2;150;155;147mQ\033[38;2;242;250;231m8\033[38;2;239;250;230m8\033[38;2;184;213;199mk\033[38;2;70;156;126mz\033[38;2;31;125;81mf\033[38;2;14;106;59m_\033[38;2;63;208;174mQ\033[38;2;70;222;200mZ\033[38;2;83;167;142mU\033[38;2;199;235;216m*\033[38;2;238;255;235mB\033[38;2;238;248;223m&\033[38;2;243;249;225m8\033[38;2;194;221;203ma\033[38;2;73;116;102mn\033[38;2;168;190;176mq\033[38;2;231;242;218mW\033[38;2;192;204;179mb\033[38;2;228;232;211mM\033[38;2;243;244;223m&\033[38;2;234;244;220mW\033[38;2;169;218;199mk\033[38;2;46;188;181mC\033[38;2;43;189;179mJ\033[38;2;136;163;159m0\033[38;2;254;253;253m \033[38;2;255;255;255m             ");
  $display("\033[38;2;255;255;255m                                     \033[38;2;254;254;254m \033[38;2;255;255;255m \033[38;2;250;250;250m@\033[38;2;227;229;227mM\033[38;2;183;192;187md\033[38;2;123;146;134mJ\033[38;2;83;121;105mu\033[38;2;61;107;92mr\033[38;2;48;106;90mj\033[38;2;47;114;97mr\033[38;2;51;120;101mr\033[38;2;54;121;101mx\033[38;2;56;120;99mx\033[38;2;56;120;98mx\033[38;2;57;120;102mx\033[38;2;57;119;102mx\033[38;2;56;119;101mx\033[38;2;56;119;102mx\033[38;2;56;123;105mx\033[38;2;62;124;108mn\033[38;2;36;66;60m+\033[38;2;6;18;15m'\033[38;2;57;105;89mj\033[38;2;52;122;104mx\033[38;2;57;119;103mx\033[38;2;47;93;81m1\033[38;2;4;14;15m'\033[38;2;15;31;30m;\033[38;2;55;85;79m1\033[38;2;15;20;23m,\033[38;2;1;0;1m \033[38;2;4;0;0m \033[38;2;11;22;21m \033[38;2;51;96;87mf\033[38;2;52;116;105mx\033[38;2;46;114;101mr\033[38;2;48;104;90mf\033[38;2;126;147;133mJ\033[38;2;236;241;223m&\033[38;2;207;212;189mh\033[38;2;199;207;184mk\033[38;2;243;249;227m8\033[38;2;210;213;198ma\033[38;2;151;156;144mQ\033[38;2;168;182;164mw\033[38;2;203;212;191mh\033[38;2;233;239;221mW\033[38;2;179;214;192mk\033[38;2;75;120;100mn\033[38;2;1;32;13m \033[38;2;8;64;37ml\033[38;2;28;96;79m?\033[38;2;19;58;47m!\033[38;2;60;95;79mf\033[38;2;199;226;205mo\033[38;2;238;251;228m8\033[38;2;185;223;199mh\033[38;2;72;131;118mv\033[38;2;117;152;138mJ\033[38;2;211;237;218m#\033[38;2;162;191;167mw\033[38;2;221;239;220mM\033[38;2;233;252;229m8\033[38;2;188;243;221m*\033[38;2;111;209;190mm\033[38;2;50;173;162mU\033[38;2;49;145;136mc\033[38;2;177;210;203mk\033[38;2;246;251;251m@\033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                                      \033[38;2;252;252;252m \033[38;2;213;212;209mo\033[38;2;146;151;146mQ\033[38;2;106;124;117mz\033[38;2;79;108;99mn\033[38;2;57;97;85mf\033[38;2;45;99;84mf\033[38;2;51;114;97mr\033[38;2;53;118;101mr\033[38;2;52;120;102mx\033[38;2;54;124;103mx\033[38;2;58;122;99mx\033[38;2;58;124;99mx\033[38;2;59;124;103mn\033[38;2;59;123;104mn\033[38;2;58;122;105mn\033[38;2;58;121;105mx\033[38;2;59;122;104mn\033[38;2;56;126;106mn\033[38;2;59;111;97mr\033[38;2;10;23;19m \033[38;2;47;89;73m?\033[38;2;57;126;106mn\033[38;2;59;120;103mx\033[38;2;50;97;84mf\033[38;2;13;24;22m,\033[38;2;3;0;1m \033[38;2;7;10;13m'\033[38;2;8;8;13m.\033[38;2;1;2;5m \033[38;2;3;2;1m \033[38;2;2;1;0m \033[38;2;9;16;15m'\033[38;2;37;68;62m+\033[38;2;53;100;89mf\033[38;2;35;70;60m+\033[38;2;71;98;84mj\033[38;2;142;157;138mL\033[38;2;233;235;214mM\033[38;2;232;236;215mM\033[38;2;206;212;189mh\033[38;2;198;203;182mb\033[38;2;198;209;191mk\033[38;2;150;169;152mO\033[38;2;197;207;188mk\033[38;2;187;197;178md\033[38;2;207;213;193ma\033[38;2;229;245;227m&\033[38;2;134;158;146mL\033[38;2;47;62;48m~\033[38;2;14;18;17m \033[38;2;6;5;4m.\033[38;2;5;10;9m.\033[38;2;53;93;85mf\033[38;2;81;133;124mc\033[38;2;46;110;98mj\033[38;2;90;138;127mz\033[38;2;157;207;193md\033[38;2;103;162;143mJ\033[38;2;156;222;208mk\033[38;2;158;238;222ma\033[38;2;97;188;174m0\033[38;2;49;131;125mu\033[38;2;28;131;125mx\033[38;2;34;201;199mL\033[38;2;48;155;153mz\033[38;2;220;217;215m*\033[38;2;255;255;255m               ");
  $display("\033[38;2;255;255;255m                                          \033[38;2;249;248;248m@\033[38;2;224;223;224mM\033[38;2;176;178;178mq\033[38;2;114;126;123mX\033[38;2;54;76;70m-\033[38;2;39;73;62m_\033[38;2;60;122;102mx\033[38;2;58;121;100mx\033[38;2;56;121;99mx\033[38;2;58;123;102mx\033[38;2;58;123;105mn\033[38;2;57;121;104mx\033[38;2;55;121;103mx\033[38;2;55;123;102mx\033[38;2;55;124;103mx\033[38;2;62;114;99mx\033[38;2;14;30;25m,\033[38;2;45;82;69m-\033[38;2;61;127;106mn\033[38;2;56;119;102mx\033[38;2;58;116;100mx\033[38;2;42;76;66m_\033[38;2;2;7;8m.\033[38;2;1;0;4m \033[38;2;0;2;5m \033[38;2;0;3;4m \033[38;2;1;3;2m \033[38;2;2;2;0m \033[38;2;0;0;0m  \033[38;2;21;33;31m;\033[38;2;46;93;83m1\033[38;2;48;109;93mj\033[38;2;57;101;85mj\033[38;2;171;192;175mq\033[38;2;159;170;150mO\033[38;2;219;228;207m*\033[38;2;238;245;225m&\033[38;2;156;165;148m0\033[38;2;163;178;159mm\033[38;2;230;246;226m&\033[38;2;118;137;123mY\033[38;2;176;187;172mq\033[38;2;159;180;169mm\033[38;2;144;158;147mQ\033[38;2;226;236;216mM\033[38;2;172;187;172mq\033[38;2;161;173;159mZ\033[38;2;183;191;177mp\033[38;2;164;174;161mm\033[38;2;159;173;158mZ\033[38;2;198;210;192mh\033[38;2;192;240;220m*\033[38;2;59;155;144mX\033[38;2;59;159;135mz\033[38;2;70;165;133mX\033[38;2;24;96;72m-\033[38;2;9;55;41ml\033[38;2;23;93;82m-\033[38;2;33;193;181mJ\033[38;2;12;255;252mw\033[38;2;47;183;183mJ\033[38;2;217;223;221m#\033[38;2;255;255;255m               ");
  $display("\033[38;2;255;255;255m                               \033[38;2;255;254;255m \033[38;2;252;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m     \033[38;2;255;254;255m \033[38;2;255;255;255m    \033[38;2;245;243;243mB\033[38;2;182;187;183mp\033[38;2;80;95;86mr\033[38;2;30;56;44mi\033[38;2;61;117;97mx\033[38;2;58;124;102mx\033[38;2;61;124;104mn\033[38;2;60;125;104mn\033[38;2;59;124;104mn\033[38;2;59;124;105mn\033[38;2;59;125;106mn\033[38;2;52;113;93mr\033[38;2;49;100;83mf\033[38;2;40;77;66m_\033[38;2;6;14;12m'\033[38;2;19;35;30m;\033[38;2;58;105;91mj\033[38;2;62;123;105mn\033[38;2;54;124;104mx\033[38;2;56;112;98mr\033[38;2;27;49;47m!\033[38;2;3;3;9m.\033[38;2;2;1;4m \033[38;2;0;3;2m \033[38;2;3;2;2m \033[38;2;2;0;1m \033[38;2;9;16;16m'\033[38;2;28;44;41ml\033[38;2;16;31;26m;\033[38;2;47;90;78m?\033[38;2;55;114;97mr\033[38;2;51;108;97mj\033[38;2;49;104;95mj\033[38;2;47;93;79m1\033[38;2;139;162;145mQ\033[38;2;180;188;173mq\033[38;2;232;235;220mW\033[38;2;185;192;173mp\033[38;2;155;173;151mO\033[38;2;138;157;142mL\033[38;2;191;217;206ma\033[38;2;65;116;109mn\033[38;2;134;155;141mL\033[38;2;217;229;210m*\033[38;2;86;126;113mv\033[38;2;167;192;177mq\033[38;2;255;255;241m@\033[38;2;249;255;235mB\033[38;2;219;235;214m#\033[38;2;158;178;162mm\033[38;2;91;125;117mc\033[38;2;48;109;99mj\033[38;2;30;97;76m?\033[38;2;18;105;87m?\033[38;2;28;133;114mx\033[38;2;41;169;150mX\033[38;2;61;188;173mC\033[38;2;90;171;172mL\033[38;2;102;201;200mm\033[38;2;155;203;201md\033[38;2;246;245;241mB\033[38;2;254;255;254m \033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                               \033[38;2;252;253;254m \033[38;2;223;248;248m8\033[38;2;197;249;244mW\033[38;2;234;252;248mB\033[38;2;255;255;254m \033[38;2;255;255;255m     \033[38;2;240;240;239m8\033[38;2;190;191;190mb\033[38;2;126;140;134mJ\033[38;2;71;104;92mr\033[38;2;51;104;85mf\033[38;2;61;121;100mx\033[38;2;37;79;68m_\033[38;2;61;114;100mx\033[38;2;56;129;107mn\033[38;2;60;126;107mn\033[38;2;61;125;108mn\033[38;2;60;124;107mnn\033[38;2;61;126;107mn\033[38;2;45;92;75m?\033[38;2;19;37;31mI\033[38;2;5;11;11m.\033[38;2;3;0;3m \033[38;2;2;0;0m \033[38;2;8;15;12m'\033[38;2;33;59;50mi\033[38;2;50;94;81m1\033[38;2;49;108;93mj\033[38;2;46;100;86mf\033[38;2;26;47;44m!\033[38;2;4;3;5m \033[38;2;2;2;2m \033[38;2;4;0;1m \033[38;2;12;23;18m \033[38;2;52;95;85mf\033[38;2;57;120;105mx\033[38;2;46;83;74m?\033[38;2;19;39;35mI\033[38;2;53;101;90mj\033[38;2;50;107;98mj\033[38;2;44;95;89mf\033[38;2;48;91;79m1\033[38;2;104;125;110mc\033[38;2;179;186;172mq\033[38;2;187;190;174mp\033[38;2;177;186;165mq\033[38;2;226;241;218mW\033[38;2;158;187;164mm\033[38;2;129;167;149mQ\033[38;2;98;128;117mz\033[38;2;233;252;235m8\033[38;2;131;166;149mQ\033[38;2;60;102;95mj\033[38;2;145;167;158m0\033[38;2;182;206;193mb\033[38;2;133;173;160m0\033[38;2;56;109;99mr\033[38;2;30;81;75m-\033[38;2;20;57;49m!\033[38;2;38;123;118mx\033[38;2;36;184;181mJ\033[38;2;66;193;187mQ\033[38;2;127;194;194mw\033[38;2;191;208;210mh\033[38;2;229;237;235m&\033[38;2;248;247;247m@\033[38;2;255;250;251m \033[38;2;255;255;255m                 ");
  $display("\033[38;2;255;255;255m                       \033[38;2;254;255;255m \033[38;2;255;255;255m    \033[38;2;254;255;255m  \033[38;2;255;255;254m \033[38;2;253;255;254m \033[38;2;253;253;253m \033[38;2;223;253;249m8\033[38;2;194;245;239mM\033[38;2;237;251;249mB\033[38;2;255;255;255m  \033[38;2;239;243;243m8\033[38;2;186;198;195mb\033[38;2;125;151;141mC\033[38;2;74;115;98mn\033[38;2;48;101;79mf\033[38;2;50;113;92mj\033[38;2;57;123;102mx\033[38;2;59;125;105mn\033[38;2;62;125;107mn\033[38;2;40;82;73m-\033[38;2;51;91;83m1\033[38;2;62;121;106mn\033[38;2;63;129;111mu\033[38;2;61;126;109mn\033[38;2;61;124;107mn\033[38;2;60;123;107mn\033[38;2;58;127;108mn\033[38;2;55;108;92mj\033[38;2;7;16;16m'\033[38;2;1;0;5m \033[38;2;2;2;5m \033[38;2;3;2;3m \033[38;2;2;0;0m \033[38;2;0;0;0m \033[38;2;4;5;6m.\033[38;2;14;27;27m,\033[38;2;21;44;40ml\033[38;2;29;43;42m!\033[38;2;10;12;14m'\033[38;2;0;0;0m  \033[38;2;29;56;47mi\033[38;2;60;117;102mx\033[38;2;50;114;102mr\033[38;2;53;116;103mr\033[38;2;26;53;47m!\033[38;2;16;31;26m;\033[38;2;86;110;98mn\033[38;2;144;163;146mQ\033[38;2;197;207;189mk\033[38;2;242;249;228m8\033[38;2;244;252;230mB\033[38;2;219;226;204m*\033[38;2;221;228;207m*\033[38;2;188;199;178md\033[38;2;163;176;155mZ\033[38;2;177;190;171mq\033[38;2;173;184;167mw\033[38;2;189;206;186mb\033[38;2;102;121;108mc\033[38;2;207;223;206mo\033[38;2;114;140;132mU\033[38;2;89;119;113mv\033[38;2;74;127;119mv\033[38;2;41;113;107mr\033[38;2;44;126;119mn\033[38;2;32;143;133mu\033[38;2;36;169;162mX\033[38;2;100;167;162mL\033[38;2;233;235;232m&\033[38;2;255;254;255m \033[38;2;255;255;255m          \033[38;2;254;255;255m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m                             \033[38;2;255;254;254m \033[38;2;253;254;253m \033[38;2;254;254;254m \033[38;2;255;254;255m \033[38;2;255;255;255m \033[38;2;252;255;255m \033[38;2;254;255;255m \033[38;2;216;226;226m#\033[38;2;125;184;176mO\033[38;2;77;174;160mJ\033[38;2;44;146;131mv\033[38;2;43;146;126mv\033[38;2;51;134;114mn\033[38;2;57;134;111mu\033[38;2;56;135;114mu\033[38;2;54;132;111mn\033[38;2;58;133;112mu\033[38;2;57;129;109mn\033[38;2;63;126;110mn\033[38;2;52;100;88mf\033[38;2;37;74;62m_\033[38;2;48;89;76m?\033[38;2;62;116;99mx\033[38;2;64;129;110mu\033[38;2;61;129;111mu\033[38;2;60;127;110mn\033[38;2;62;130;111mu\033[38;2;36;71;64m_\033[38;2;0;2;6m \033[38;2;1;2;4m \033[38;2;1;3;2m   \033[38;2;2;1;0m \033[38;2;0;0;4m \033[38;2;0;0;0m \033[38;2;8;11;9m.\033[38;2;38;55;54m~\033[38;2;24;42;36ml\033[38;2;16;26;22m,\033[38;2;30;54;50mi\033[38;2;58;113;102mx\033[38;2;51;113;102mr\033[38;2;52;114;102mr\033[38;2;37;71;61m+\033[38;2;1;4;1m \033[38;2;62;69;59m-\033[38;2;213;224;204mo\033[38;2;254;255;241m@\033[38;2;246;254;231mB\033[38;2;242;251;227m8\033[38;2;243;253;229m8\033[38;2;242;252;228m8\033[38;2;238;245;222m&\033[38;2;241;244;222m&\033[38;2;181;189;168mq\033[38;2;157;172;155mO\033[38;2;139;152;137mC\033[38;2;150;160;146m0\033[38;2;161;179;158mm\033[38;2;117;145;133mU\033[38;2;172;189;175mq\033[38;2;109;150;134mU\033[38;2;121;168;159mQ\033[38;2;113;181;171m0\033[38;2;35;158;149mz\033[38;2;45;173;167mU\033[38;2;187;223;221mo\033[38;2;255;255;255m                       ");
  $display("\033[38;2;255;255;255m                      \033[38;2;254;255;254m \033[38;2;227;235;234mW\033[38;2;213;229;226m#\033[38;2;234;241;239m8\033[38;2;207;237;237mM\033[38;2;157;234;233ma\033[38;2;178;244;244m#\033[38;2;226;253;252mB\033[38;2;250;254;255m \033[38;2;255;254;255m \033[38;2;255;254;254m \033[38;2;255;255;255m \033[38;2;245;241;240mB\033[38;2;152;155;151m0\033[38;2;63;91;80mf\033[38;2;44;116;94mj\033[38;2;51;128;107mn\033[38;2;51;125;104mx\033[38;2;46;122;99mr\033[38;2;54;118;99mr\033[38;2;52;122;102mx\033[38;2;52;129;110mn\033[38;2;51;134;114mn\033[38;2;55;137;117mu\033[38;2;55;128;110mn\033[38;2;61;130;110mu\033[38;2;65;132;111mu\033[38;2;61;121;100mx\033[38;2;38;84;66m-\033[38;2;28;57;44mi\033[38;2;34;67;54m~\033[38;2;48;93;78m1\033[38;2;55;109;93mj\033[38;2;57;115;100mr\033[38;2;63;110;98mr\033[38;2;25;37;37mI\033[38;2;1;2;4m \033[38;2;1;3;2m \033[38;2;1;3;3m  \033[38;2;2;2;2m \033[38;2;1;1;6m \033[38;2;0;0;2m \033[38;2;10;23;18m \033[38;2;65;113;103mx\033[38;2;58;123;104mn\033[38;2;57;117;99mx\033[38;2;52;109;96mj\033[38;2;52;114;104mr\033[38;2;52;113;105mr\033[38;2;51;112;102mr\033[38;2;34;67;60m+\033[38;2;3;5;4m \033[38;2;0;0;0m \033[38;2;33;38;34ml\033[38;2;142;160;146mQ\033[38;2;231;249;226m&\033[38;2;246;255;233mB\033[38;2;245;251;228m8\033[38;2;244;249;227m8\033[38;2;241;251;228m8\033[38;2;243;251;227m8\033[38;2;226;237;214mM\033[38;2;155;172;153mO\033[38;2;115;154;142mJ\033[38;2;48;103;92mj\033[38;2;132;163;152mQ\033[38;2;102;133;128mX\033[38;2;93;129;118mc\033[38;2;127;194;178mm\033[38;2;79;173;165mC\033[38;2;57;178;170mJ\033[38;2;71;144;137mz\033[38;2;172;194;188mp\033[38;2;249;252;253m@\033[38;2;252;254;252m \033[38;2;255;255;255m          \033[38;2;253;253;252m \033[38;2;245;249;245mB\033[38;2;238;247;242mB\033[38;2;233;248;246mB\033[38;2;244;252;252m@\033[38;2;255;255;255m  \033[38;2;254;255;255m \033[38;2;255;255;255m    ");
  $display("\033[38;2;255;255;255m        \033[38;2;254;254;253m \033[38;2;254;254;252m \033[38;2;246;253;252m@\033[38;2;233;251;251mB\033[38;2;249;254;254m \033[38;2;255;255;255m \033[38;2;255;255;254m \033[38;2;254;254;254m \033[38;2;255;255;255m     \033[38;2;202;204;201mh\033[38;2;105;137;125mX\033[38;2;63;125;112mu\033[38;2;46;124;114mx\033[38;2;49;127;110mn\033[38;2;37;139;123mn\033[38;2;34;172;165mX\033[38;2;37;196;191mC\033[38;2;85;224;222mq\033[38;2;148;245;241mo\033[38;2;212;254;254m8\033[38;2;224;251;248m8\033[38;2;173;226;223ma\033[38;2;63;130;118mu\033[38;2;29;90;73m-\033[38;2;56;108;93mj\033[38;2;62;108;91mr\033[38;2;86;112;99mn\033[38;2;116;135;126mY\033[38;2;139;160;148mQ\033[38;2;156;176;164mZ\033[38;2;139;161;152mQ\033[38;2;114;140;129mY\033[38;2;95;126;114mc\033[38;2;77;114;102mn\033[38;2;65;104;92mr\033[38;2;58;101;86mj\033[38;2;50;95;79m1\033[38;2;45;95;77m1\033[38;2;41;95;76m?\033[38;2;38;82;67m-\033[38;2;28;49;42m!\033[38;2;18;27;24m,\033[38;2;11;20;17m \033[38;2;9;18;15m'\033[38;2;12;20;18m \033[38;2;12;13;13m'\033[38;2;3;3;3m \033[38;2;1;3;2m   \033[38;2;2;2;4m \033[38;2;1;2;6m \033[38;2;1;0;2m \033[38;2;8;22;17m \033[38;2;58;110;94mr\033[38;2;54;119;102mx\033[38;2;54;118;102mx\033[38;2;54;117;103mx\033[38;2;53;115;103mr\033[38;2;52;113;102mr\033[38;2;52;112;99mr\033[38;2;30;59;54mi\033[38;2;1;2;4m \033[38;2;2;1;3m \033[38;2;0;0;0m \033[38;2;4;11;6m.\033[38;2;76;96;84mj\033[38;2;185;208;189mb\033[38;2;236;252;229m8\033[38;2;249;254;233mB\033[38;2;245;249;229m8\033[38;2;243;248;224m8\033[38;2;241;250;225m8\033[38;2;230;247;225m&\033[38;2;111;167;153mL\033[38;2;29;116;107mj\033[38;2;32;109;100mf\033[38;2;30;115;106mj\033[38;2;46;157;143mz\033[38;2;56;223;216mZ\033[38;2;31;191;194mC\033[38;2;102;179;173mQ\033[38;2;228;235;233mW\033[38;2;255;255;255m  \033[38;2;254;254;255m \033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;235;251;247mB\033[38;2;165;232;220ma\033[38;2;122;223;202mp\033[38;2;113;215;191mw\033[38;2;105;216;186mm\033[38;2;106;221;200mw\033[38;2;136;223;203md\033[38;2;236;248;241m8\033[38;2;255;255;255m \033[38;2;252;255;255m \033[38;2;253;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m        \033[38;2;253;255;254m \033[38;2;254;254;252m \033[38;2;219;249;247m8\033[38;2;113;234;221md\033[38;2;118;238;232mk\033[38;2;192;251;252mW\033[38;2;242;254;254m@\033[38;2;255;254;253m \033[38;2;255;255;255m   \033[38;2;230;230;228mW\033[38;2;130;149;140mC\033[38;2;44;92;79m?\033[38;2;37;97;82m1\033[38;2;50;109;92mj\033[38;2;91;130;124mz\033[38;2;139;168;159m0\033[38;2;185;205;197mk\033[38;2;224;234;232mW\033[38;2;227;244;240m&\033[38;2;222;249;248m8\033[38;2;186;248;244mM\033[38;2;116;239;232mk\033[38;2;124;248;242ma\033[38;2;72;222;217mm\033[38;2;43;202;194mL\033[38;2;91;198;189mO\033[38;2;164;208;202mb\033[38;2;223;232;219mM\033[38;2;250;252;240m@\033[38;2;255;255;252m \033[38;2;255;255;251m  \033[38;2;255;255;252m \033[38;2;255;255;248m \033[38;2;255;255;242m@\033[38;2;245;246;233m8\033[38;2;227;229;216mM\033[38;2;216;216;203mo\033[38;2;194;196;185mb\033[38;2;163;167;159mZ\033[38;2;129;136;128mU\033[38;2;93;101;92mn\033[38;2;67;73;68m?\033[38;2;43;47;46mi\033[38;2;21;24;24m,\033[38;2;7;6;6m.\033[38;2;0;0;0m    \033[38;2;0;2;1m \033[38;2;1;3;2m \033[38;2;1;2;3m \033[38;2;1;2;6m \033[38;2;4;0;4m \033[38;2;6;13;10m.\033[38;2;55;102;89mj\033[38;2;56;119;104mx\033[38;2;55;117;104mx\033[38;2;55;117;106mx\033[38;2;54;114;104mr\033[38;2;55;113;102mr\033[38;2;52;109;96mj\033[38;2;23;49;45m!\033[38;2;2;1;4m \033[38;2;1;2;3m \033[38;2;1;3;2m \033[38;2;1;0;0m \033[38;2;0;0;0m \033[38;2;22;34;31mI\033[38;2;96;121;108mv\033[38;2;176;204;182md\033[38;2;227;247;224mW\033[38;2;244;255;231mB\033[38;2;248;253;230mB\033[38;2;240;249;229m8\033[38;2;120;169;155mQ\033[38;2;29;117;108mj\033[38;2;29;120;110mr\033[38;2;23;131;123mx\033[38;2;21;187;182mU\033[38;2;16;251;253mw\033[38;2;55;202;198mQ\033[38;2;212;225;222m#\033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m       \033[38;2;254;254;255m \033[38;2;162;242;238m*\033[38;2;57;231;222mm\033[38;2;84;237;229mp\033[38;2;106;239;228mb\033[38;2;77;234;224mq\033[38;2;79;223;204mm\033[38;2;101;210;177mZ\033[38;2;171;214;192mb\033[38;2;246;251;246m@\033[38;2;255;254;255m \033[38;2;253;255;254m \033[38;2;255;255;253m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m        \033[38;2;254;255;254m \033[38;2;254;255;253m \033[38;2;255;255;255m \033[38;2;227;248;247m8\033[38;2;125;229;219mb\033[38;2;91;234;224mp\033[38;2;160;251;245m*\033[38;2;244;251;254m@\033[38;2;255;255;255m \033[38;2;246;244;244mB\033[38;2;162;171;162mZ\033[38;2;62;101;84mj\033[38;2;53;104;87mj\033[38;2;96;142;127mX\033[38;2;158;182;172mm\033[38;2;217;224;218m#\033[38;2;255;254;253m \033[38;2;255;255;255m \033[38;2;251;247;247m@\033[38;2;237;232;233m&\033[38;2;221;217;215m*\033[38;2;191;193;189mb\033[38;2;117;163;155mL\033[38;2;60;186;179mC\033[38;2;64;223;215mm\033[38;2;113;244;243mh\033[38;2;135;254;250mo\033[38;2;108;247;243mk\033[38;2;101;237;234mb\033[38;2;133;214;200mp\033[38;2;150;185;173mm\033[38;2;162;178;163mm\033[38;2;168;168;160mZ\033[38;2;173;175;168mw\033[38;2;180;183;175mq\033[38;2;190;191;180md\033[38;2;201;202;190mk\033[38;2;209;211;199ma\033[38;2;220;221;210m*\033[38;2;233;234;222mW\033[38;2;243;244;231m8\033[38;2;252;254;240m@\033[38;2;255;255;245m@@\033[38;2;255;255;242m@\033[38;2;242;242;230m8\033[38;2;221;220;210m*\033[38;2;187;187;180mp\033[38;2;147;148;140mL\033[38;2;105;105;98mu\033[38;2;58;59;54m_\033[38;2;20;21;20m,\033[38;2;0;0;1m \033[38;2;0;0;0m    \033[38;2;0;0;1m \033[38;2;43;78;69m-\033[38;2;56;122;104mx\033[38;2;53;117;103mx\033[38;2;54;113;105mr\033[38;2;50;115;106mr\033[38;2;54;114;102mr\033[38;2;54;110;94mr\033[38;2;25;50;44m!\033[38;2;1;1;6m  \033[38;2;1;2;5m \033[38;2;2;2;3m \033[38;2;2;2;2m \033[38;2;0;0;0m \033[38;2;0;1;2m \033[38;2;19;34;32m;\033[38;2;66;105;96mr\033[38;2;130;185;167mO\033[38;2;187;234;213mo\033[38;2;185;231;208ma\033[38;2;88;159;144mU\033[38;2;29;117;110mj\033[38;2;32;122;114mr\033[38;2;23;135;132mn\033[38;2;24;206;204mL\033[38;2;25;240;237mm\033[38;2;112;185;182mO\033[38;2;254;252;251m \033[38;2;255;255;255m     \033[38;2;254;255;255m  \033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;255;255;253m \033[38;2;229;252;252mB\033[38;2;136;245;241ma\033[38;2;96;243;235mb\033[38;2;158;249;246m*\033[38;2;223;252;253mB\033[38;2;232;255;255m@\033[38;2;132;246;248ma\033[38;2;68;231;226mw\033[38;2;84;221;195mm\033[38;2;121;202;169mZ\033[38;2;223;237;226mW\033[38;2;255;255;255m \033[38;2;254;254;255m \033[38;2;254;255;254m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m           \033[38;2;255;255;254m \033[38;2;248;254;252m@\033[38;2;172;236;230mo\033[38;2;107;234;224md\033[38;2;154;249;247m*\033[38;2;182;236;231m*\033[38;2;98;152;141mU\033[38;2;89;125;112mv\033[38;2;165;182;174mw\033[38;2;227;234;230mW\033[38;2;255;255;255m \033[38;2;235;232;231mW\033[38;2;171;172;170mw\033[38;2;122;130;128mY\033[38;2;89;107;101mn\033[38;2;71;98;89mr\033[38;2;57;90;82mf\033[38;2;41;86;73m-\033[38;2;37;92;74m?\033[38;2;31;112;86mf\033[38;2;35;163;132mc\033[38;2;35;212;188mL\033[38;2;33;236;218mZ\033[38;2;81;243;233md\033[38;2;120;246;242mh\033[38;2;87;239;233md\033[38;2;23;213;201mL\033[38;2;18;153;137mu\033[38;2;17;91;72m_\033[38;2;4;38;27m,\033[38;2;4;24;14m'\033[38;2;9;25;18m \033[38;2;7;25;17m \033[38;2;10;24;18m \033[38;2;14;22;17m \033[38;2;19;24;21m,\033[38;2;25;34;29mI\033[38;2;35;42;36ml\033[38;2;48;52;45m~\033[38;2;62;64;57m_\033[38;2;75;80;71m1\033[38;2;98;102;93mn\033[38;2;123;128;119mX\033[38;2;149;154;146mQ\033[38;2;178;184;175mq\033[38;2;210;213;202ma\033[38;2;234;234;222mW\033[38;2;240;241;226m&\033[38;2;223;225;210m#\033[38;2;191;193;181md\033[38;2;146;148;139mL\033[38;2;90;89;82mr\033[38;2;40;45;37m!\033[38;2;24;33;28m;\033[38;2;23;41;37mI\033[38;2;36;80;68m_\033[38;2;53;120;101mx\033[38;2;54;119;104mx\033[38;2;55;114;106mx\033[38;2;49;116;105mr\033[38;2;53;115;105mx\033[38;2;49;107;96mj\033[38;2;31;62;56m~\033[38;2;5;8;11m.\033[38;2;1;1;6m \033[38;2;1;2;6m \033[38;2;1;2;4m \033[38;2;1;1;1m \033[38;2;3;3;4m \033[38;2;8;7;11m.\033[38;2;3;0;5m \033[38;2;0;3;4m \033[38;2;5;27;27m,\033[38;2;29;69;72m+\033[38;2;40;122;116mx\033[38;2;38;149;138mv\033[38;2;34;154;148mc\033[38;2;32;154;142mv\033[38;2;16;157;148mv\033[38;2;16;220;212mQ\033[38;2;40;219;215mO\033[38;2;172;204;203mb\033[38;2;255;255;255m        \033[38;2;243;252;250m@\033[38;2;204;247;243mW\033[38;2;138;240;233mh\033[38;2;96;242;234mb\033[38;2;135;246;246mo\033[38;2;192;253;251mW\033[38;2;220;247;247m8\033[38;2;247;253;252m@\033[38;2;220;254;253mB\033[38;2;98;242;239mb\033[38;2;60;236;229mw\033[38;2;77;225;203mm\033[38;2;116;206;176mm\033[38;2;224;239;228mW\033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;254;255;254m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m            \033[38;2;255;255;253m \033[38;2;255;254;254m \033[38;2;194;244;240mM\033[38;2;116;235;228mb\033[38;2;118;236;226mb\033[38;2;202;231;226m#\033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;208;202;202ma\033[38;2;109;110;109mv\033[38;2;42;62;54m~\033[38;2;34;72;63m+\033[38;2;41;99;87m1\033[38;2;47;111;95mj\033[38;2;47;130;105mx\033[38;2;48;155;120mv\033[38;2;53;177;134mX\033[38;2;59;196;147mJ\033[38;2;54;191;138mY\033[38;2;50;183;132mX\033[38;2;46;169;131mz\033[38;2;33;163;142mc\033[38;2;24;193;181mU\033[38;2;40;221;213mO\033[38;2;99;244;240mb\033[38;2;107;245;245mk\033[38;2;55;221;215mZ\033[38;2;26;189;176mU\033[38;2;33;157;139mv\033[38;2;39;128;108mx\033[38;2;40;110;93mj\033[38;2;38;99;80m1\033[38;2;35;89;71m-\033[38;2;32;77;63m_\033[38;2;30;68;56m~\033[38;2;20;49;42ml\033[38;2;11;32;25m,\033[38;2;5;15;10m'\033[38;2;0;2;0m \033[38;2;0;0;0m    \033[38;2;2;9;7m.\033[38;2;11;17;14m'\033[38;2;31;35;31mI\033[38;2;56;62;56m_\033[38;2;85;93;83mr\033[38;2;140;146;133mC\033[38;2;215;221;205mo\033[38;2;251;255;237m@\033[38;2;247;252;231mB\033[38;2;215;224;205m*\033[38;2;165;184;166mw\033[38;2;118;150;132mJ\033[38;2;79;126;107mu\033[38;2;50;108;92mj\033[38;2;50;111;100mr\033[38;2;53;114;103mr\033[38;2;51;112;104mr\033[38;2;47;106;98mj\033[38;2;38;82;72m-\033[38;2;20;36;34mI\033[38;2;1;1;5m \033[38;2;3;0;4m \033[38;2;2;2;3m \033[38;2;2;1;1m \033[38;2;3;4;4m \033[38;2;18;33;31m;\033[38;2;12;22;23m,\033[38;2;1;2;3m \033[38;2;0;1;1m \033[38;2;0;1;2m \033[38;2;4;15;13m'\033[38;2;14;38;38mI\033[38;2;17;64;64m~\033[38;2;28;105;101mf\033[38;2;51;168;158mY\033[38;2;50;205;197mQ\033[38;2;65;181;181mC\033[38;2;214;225;220m#\033[38;2;255;255;255m   \033[38;2;255;255;254m \033[38;2;249;252;251m@\033[38;2;230;248;245m8\033[38;2;198;243;237mM\033[38;2;156;238;230ma\033[38;2;115;234;221mb\033[38;2;91;238;226md\033[38;2;98;238;234mb\033[38;2;109;244;238mk\033[38;2;123;247;241mh\033[38;2;107;243;243mk\033[38;2;162;247;248m#\033[38;2;240;253;254m@\033[38;2;165;249;247m#\033[38;2;63;241;232mq\033[38;2;63;234;224mw\033[38;2;88;218;193mm\033[38;2;141;211;183mq\033[38;2;244;250;243mB\033[38;2;255;254;255m \033[38;2;252;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m           \033[38;2;255;254;255m \033[38;2;255;254;254m \033[38;2;255;255;252m \033[38;2;255;255;255m \033[38;2;201;241;239mM\033[38;2;129;237;227mk\033[38;2;208;255;255m8\033[38;2;198;221;219mo\033[38;2;95;110;102mu\033[38;2;30;53;44m!\033[38;2;33;81;69m_\033[38;2;49;109;99mj\033[38;2;51;115;105mr\033[38;2;53;112;101mr\033[38;2;43;133;106mx\033[38;2;60;190;142mU\033[38;2;52;170;125mz\033[38;2;51;148;111mu\033[38;2;48;126;97mr\033[38;2;48;114;89mj\033[38;2;54;121;101mx\033[38;2;58;129;108mn\033[38;2;55;139;116mu\033[38;2;47;156;134mc\033[38;2;38;179;163mY\033[38;2;36;208;195mL\033[38;2;68;234;228mq\033[38;2;101;248;244mk\033[38;2;82;244;237md\033[38;2;66;237;232mq\033[38;2;53;220;211mO\033[38;2;44;198;181mC\033[38;2;41;166;149mz\033[38;2;30;122;108mr\033[38;2;26;76;66m+\033[38;2;20;43;37mI\033[38;2;15;28;26m,\033[38;2;10;21;20m \033[38;2;9;19;16m'\033[38;2;9;18;15m'\033[38;2;9;18;14m'\033[38;2;8;17;14m'\033[38;2;6;15;12m'\033[38;2;5;15;11m'\033[38;2;5;15;12m'\033[38;2;3;13;10m.\033[38;2;3;12;9m.\033[38;2;0;8;5m \033[38;2;0;0;0m \033[38;2;0;2;0m \033[38;2;18;22;19m,\033[38;2;70;75;68m?\033[38;2;135;144;132mJ\033[38;2;217;224;209m*\033[38;2;255;255;246m \033[38;2;255;255;243m@\033[38;2;238;241;224m&\033[38;2;169;184;171mw\033[38;2;72;110;95mx\033[38;2;47;100;86mf\033[38;2;52;114;102mr\033[38;2;47;111;102mr\033[38;2;38;92;82m?\033[38;2;34;74;65m_\033[38;2;15;33;31m;\033[38;2;3;5;6m \033[38;2;1;1;1m \033[38;2;2;3;2m \033[38;2;4;1;2m \033[38;2;24;44;40ml\033[38;2;29;67;58m~\033[38;2;18;38;36mI\033[38;2;7;10;9m.\033[38;2;3;14;12m.\033[38;2;43;83;79m?\033[38;2;30;55;54mi\033[38;2;5;9;12m.\033[38;2;11;18;15m'\033[38;2;161;160;158mO\033[38;2;234;236;236m&\033[38;2;225;227;228mM\033[38;2;252;252;247m@\033[38;2;250;253;252m@\033[38;2;226;248;241m8\033[38;2;195;243;232mM\033[38;2;160;236;226ma\033[38;2;138;233;226mk\033[38;2;125;232;223mb\033[38;2;135;237;225mk\033[38;2;162;241;234mo\033[38;2;188;243;241mM\033[38;2;197;247;242mW\033[38;2;194;247;241mM\033[38;2;201;248;244mW\033[38;2;213;252;248m&\033[38;2;188;246;247mM\033[38;2;192;251;248mW\033[38;2;217;254;252m8\033[38;2;106;241;239mk\033[38;2;55;238;229mw\033[38;2;76;227;207mm\033[38;2;106;210;177mZ\033[38;2;205;232;217m*\033[38;2;255;255;254m \033[38;2;254;254;253m \033[38;2;253;255;254m \033[38;2;255;255;255m   ");
  $display("\033[38;2;255;255;255m           \033[38;2;254;254;255m  \033[38;2;253;254;255m \033[38;2;255;255;255m \033[38;2;242;255;254m@\033[38;2;124;237;227mk\033[38;2;75;222;217mw\033[38;2;30;134;126mn\033[38;2;30;98;88m1\033[38;2;51;109;100mr\033[38;2;51;113;102mr\033[38;2;48;111;98mj\033[38;2;49;111;101mr\033[38;2;46;108;94mj\033[38;2;50;167;125mz\033[38;2;49;153;115mv\033[38;2;45;100;83mf\033[38;2;57;121;103mx\033[38;2;57;129;110mn\033[38;2;57;132;113mu\033[38;2;56;134;114mu\033[38;2;60;134;114mu\033[38;2;61;134;114mu\033[38;2;58;136;116mu\033[38;2;55;140;122mv\033[38;2;45;157;136mc\033[38;2;41;176;160mY\033[38;2;47;196;185mC\033[38;2;56;206;197m0\033[38;2;51;198;192mQ\033[38;2;57;210;206mO\033[38;2;67;226;223mw\033[38;2;61;221;219mm\033[38;2;44;190;188mC\033[38;2;27;144;143mu\033[38;2;25;117;114mj\033[38;2;37;117;107mr\033[38;2;47;116;101mr\033[38;2;58;115;99mr\033[38;2;57;117;100mx\033[38;2;55;115;98mrr\033[38;2;55;114;96mr\033[38;2;52;110;92mj\033[38;2;50;103;88mf\033[38;2;46;94;81m1\033[38;2;39;84;72m-\033[38;2;32;70;59m+\033[38;2;22;49;39ml\033[38;2;10;26;20m \033[38;2;3;11;7m.\033[38;2;0;3;2m \033[38;2;0;4;3m \033[38;2;29;40;34ml\033[38;2;85;97;87mr\033[38;2;173;185;169mw\033[38;2;244;250;230m8\033[38;2;255;255;246m \033[38;2;227;231;215mM\033[38;2;123;138;125mU\033[38;2;49;86;76m?\033[38;2;43;104;93mf\033[38;2;46;111;99mj\033[38;2;42;98;87m1\033[38;2;31;72;65m+\033[38;2;26;47;43m!\033[38;2;9;16;14m'\033[38;2;0;2;0m \033[38;2;4;0;1m \033[38;2;4;11;11m.\033[38;2;31;63;57m~\033[38;2;35;71;65m_\033[38;2;17;47;41ml\033[38;2;19;96;93m?\033[38;2;65;198;190mQ\033[38;2;29;87;85m?\033[38;2;6;27;26m,\033[38;2;36;97;89m1\033[38;2;141;164;161m0\033[38;2;245;255;255m@\033[38;2;221;250;246m8\033[38;2;188;241;235m#\033[38;2;152;239;223ma\033[38;2;144;235;221mh\033[38;2;155;238;229ma\033[38;2;188;244;238mM\033[38;2;220;249;245m8\033[38;2;238;252;251m@\033[38;2;252;254;254m \033[38;2;255;255;255m     \033[38;2;255;255;253m \033[38;2;242;254;252m@\033[38;2;224;254;251mB\033[38;2;168;249;247m#\033[38;2;65;237;229mq\033[38;2;67;230;210mm\033[38;2;100;212;181mZ\033[38;2;180;224;203mh\033[38;2;254;254;251m \033[38;2;254;255;255m \033[38;2;254;255;254m \033[38;2;255;254;254m \033[38;2;255;255;255m   ");
  $display("\033[38;2;255;255;255m             \033[38;2;255;255;253m \033[38;2;249;255;253m \033[38;2;166;220;210mk\033[38;2;64;173;168mJ\033[38;2;32;146;143mv\033[38;2;39;126;114mx\033[38;2;46;114;103mr\033[38;2;48;110;100mr\033[38;2;49;111;100mr\033[38;2;50;111;101mr\033[38;2;51;113;102mr\033[38;2;50;112;95mj\033[38;2;43;132;100mx\033[38;2;50;136;106mn\033[38;2;52;117;98mr\033[38;2;52;122;103mx\033[38;2;52;127;106mn\033[38;2;57;129;109mn\033[38;2;57;130;109mn\033[38;2;57;130;110mn\033[38;2;59;132;112mu\033[38;2;61;134;114mu\033[38;2;64;133;114mu\033[38;2;60;133;114mu\033[38;2;59;137;117mu\033[38;2;55;131;113mn\033[38;2;15;70;59m~\033[38;2;0;37;36m;\033[38;2;3;50;51ml\033[38;2;8;86;81m_\033[38;2;29;149;138mv\033[38;2;52;205;195mQ\033[38;2;59;229;223mm\033[38;2;75;238;234mp\033[38;2;76;235;227mq\033[38;2;56;203;189mQ\033[38;2;50;153;139mz\033[38;2;55;139;122mv\033[38;2;57;137;121mv\033[38;2;62;130;115mu\033[38;2;66;129;112mu\033[38;2;63;130;111mu\033[38;2;59;132;112mu\033[38;2;60;129;111mu\033[38;2;62;130;112mu\033[38;2;63;129;111mu\033[38;2;60;125;107mn\033[38;2;50;106;89mj\033[38;2;29;70;56m~\033[38;2;8;31;21m,\033[38;2;1;10;5m.\033[38;2;0;4;3m \033[38;2;0;0;0m \033[38;2;3;8;9m.\033[38;2;61;74;66m?\033[38;2;162;180;162mm\033[38;2;234;246;228m&\033[38;2;255;255;243m@\033[38;2;205;209;193mh\033[38;2;103;120;107mc\033[38;2;41;81;68m-\033[38;2;32;83;71m-\033[38;2;40;91;79m?\033[38;2;38;81;70m-\033[38;2;32;60;53m~\033[38;2;16;29;25m,\033[38;2;4;6;6m.\033[38;2;1;0;4m \033[38;2;6;13;15m'\033[38;2;24;55;51mi\033[38;2;22;77;72m_\033[38;2;46;180;171mU\033[38;2;38;153;149mc\033[38;2;5;29;25m,\033[38;2;0;16;11m.\033[38;2;45;142;139mv\033[38;2;54;143;137mc\033[38;2;156;218;211mk\033[38;2;193;250;243mW\033[38;2;213;251;246m&\033[38;2;238;255;253m@\033[38;2;255;255;255m           \033[38;2;255;254;254m \033[38;2;247;254;254m@\033[38;2;221;253;253mB\033[38;2;136;246;239ma\033[38;2;61;236;222mw\033[38;2;85;217;195mZ\033[38;2;157;215;195md\033[38;2;249;253;250m@\033[38;2;255;254;255m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m        \033[38;2;255;255;254m \033[38;2;255;255;255m   \033[38;2;254;253;255m \033[38;2;227;247;244m8\033[38;2;118;197;186mm\033[38;2;31;121;109mr\033[38;2;35;98;90m1\033[38;2;44;105;97mj\033[38;2;44;108;95mj\033[38;2;46;107;96mj\033[38;2;46;110;98mj\033[38;2;47;111;101mr\033[38;2;50;111;103mr\033[38;2;51;112;103mr\033[38;2;53;113;102mr\033[38;2;43;106;92mf\033[38;2;43;110;92mj\033[38;2;53;121;104mx\033[38;2;52;122;106mx\033[38;2;52;124;104mx\033[38;2;54;125;105mx\033[38;2;56;126;106mn\033[38;2;58;127;107mnn\033[38;2;59;128;108mn\033[38;2;60;130;107mn\033[38;2;57;132;107mn\033[38;2;63;132;110mu\033[38;2;44;96;79m1\033[38;2;10;33;25m,\033[38;2;4;11;8m.\033[38;2;10;23;19m \033[38;2;39;79;66m_\033[38;2;55;127;104mn\033[38;2;55;136;119mu\033[38;2;47;149;135mc\033[38;2;45;167;151mX\033[38;2;52;179;165mU\033[38;2;51;176;165mU\033[38;2;40;173;163mY\033[38;2;60;209;197m0\033[38;2;63;205;196m0\033[38;2;46;168;156mX\033[38;2;48;138;120mu\033[38;2;58;125;104mn\033[38;2;62;127;107mn\033[38;2;60;128;106mn\033[38;2;61;127;108mn\033[38;2;62;125;109mn\033[38;2;61;125;108mn\033[38;2;59;125;107mn\033[38;2;57;117;101mx\033[38;2;41;90;77m?\033[38;2;18;49;41ml\033[38;2;8;18;16m'\033[38;2;3;9;6m.\033[38;2;0;8;6m \033[38;2;0;1;0m \033[38;2;3;12;7m.\033[38;2;60;85;75m1\033[38;2;148;185;171mm\033[38;2;208;237;221m#\033[38;2;240;248;236m8\033[38;2;203;206;200mh\033[38;2;120;130;125mY\033[38;2;60;74;68m?\033[38;2;24;41;35mI\033[38;2;18;36;30m;\033[38;2;12;32;25m,\033[38;2;1;13;9m.\033[38;2;0;0;0m \033[38;2;1;0;1m \033[38;2;13;16;14m'\033[38;2;27;53;49mi\033[38;2;49;92;90mf\033[38;2;28;54;49mi\033[38;2;11;25;23m,\033[38;2;0;10;7m.\033[38;2;30;90;87m?\033[38;2;46;121;113mx\033[38;2;87;100;98mn\033[38;2;179;193;192md\033[38;2;185;205;202mk\033[38;2;194;211;210ma\033[38;2;210;221;221m*\033[38;2;221;227;225mM\033[38;2;234;234;232m&\033[38;2;249;243;244mB\033[38;2;255;253;252m \033[38;2;255;255;255m  \033[38;2;253;255;254m \033[38;2;254;254;255m  \033[38;2;255;255;255m \033[38;2;236;253;250mB\033[38;2;218;249;248m8\033[38;2;204;251;252m&\033[38;2;122;244;236mh\033[38;2;68;225;205mm\033[38;2;143;219;202md\033[38;2;238;246;240m8\033[38;2;255;255;253m \033[38;2;254;255;255m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m        \033[38;2;253;252;251m \033[38;2;236;234;229m&\033[38;2;231;231;226mW\033[38;2;248;249;246m@\033[38;2;237;249;244mB\033[38;2;158;213;199mb\033[38;2;85;143;134mX\033[38;2;66;106;103mx\033[38;2;50;93;82m1\033[38;2;39;88;77m?\033[38;2;38;94;83m?\033[38;2;42;101;90mf\033[38;2;45;107;96mj\033[38;2;47;112;100mr\033[38;2;51;111;100mr\033[38;2;51;110;101mr\033[38;2;50;112;101mr\033[38;2;50;112;99mr\033[38;2;50;111;96mj\033[38;2;53;117;105mx\033[38;2;53;118;108mx\033[38;2;55;121;105mx\033[38;2;56;123;103mx\033[38;2;58;123;103mx\033[38;2;59;123;103mn\033[38;2;59;124;104mnn\033[38;2;59;127;104mn\033[38;2;58;130;105mn\033[38;2;57;121;99mx\033[38;2;32;79;63m_\033[38;2;13;41;30m;\033[38;2;23;53;41m!\033[38;2;62;110;95mr\033[38;2;65;134;113mu\033[38;2;60;130;111mu\033[38;2;64;126;110muu\033[38;2;59;127;109mn\033[38;2;57;126;105mn\033[38;2;54;128;105mn\033[38;2;47;147;128mv\033[38;2;52;187;175mC\033[38;2;67;229;221mw\033[38;2;70;236;231mq\033[38;2;55;207;196m0\033[38;2;43;169;153mX\033[38;2;47;139;123mu\033[38;2;57;124;105mn\033[38;2;60;123;100mx\033[38;2;56;125;102mx\033[38;2;58;124;104mn\033[38;2;60;124;106mn\033[38;2;62;124;108mn\033[38;2;56;117;102mx\033[38;2;47;99;85mf\033[38;2;28;62;52mi\033[38;2;11;29;22m,\033[38;2;4;16;11m'\033[38;2;4;11;9m.\033[38;2;4;7;6m.\033[38;2;0;4;2m \033[38;2;9;28;23m,\033[38;2;48;93;76m1\033[38;2;77;147;117mc\033[38;2;104;160;136mJ\033[38;2;138;173;158m0\033[38;2;151;175;164mZ\033[38;2;134;149;141mC\033[38;2;105;119;111mc\033[38;2;95;113;106mu\033[38;2;85;111;101mn\033[38;2;104;129;114mz\033[38;2;155;170;156mO\033[38;2;192;201;186mb\033[38;2;208;213;199ma\033[38;2;211;218;201mo\033[38;2;208;225;205mo\033[38;2;160;202;185mp\033[38;2;81;151;135mX\033[38;2;30;98;87m?\033[38;2;30;80;70m_\033[38;2;24;56;46m!\033[38;2;25;69;58m~\033[38;2;33;106;93mf\033[38;2;40;120;113mx\033[38;2;46;142;135mv\033[38;2;49;156;152mX\033[38;2;61;168;162mU\033[38;2;79;181;170mL\033[38;2;107;188;182mO\033[38;2;189;218;219ma\033[38;2;253;254;252m \033[38;2;253;254;254m  \033[38;2;255;255;253m \033[38;2;190;243;241mM\033[38;2;116;237;234mk\033[38;2;154;247;244m*\033[38;2;121;242;233mk\033[38;2;88;227;216mq\033[38;2;159;227;215mh\033[38;2;242;251;249m@\033[38;2;255;255;255m \033[38;2;254;255;253m \033[38;2;255;254;254m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m        \033[38;2;254;253;253m \033[38;2;232;230;224mW\033[38;2;167;170;160mZ\033[38;2;117;132;122mX\033[38;2;118;140;130mU\033[38;2;153;172;168mZ\033[38;2;185;198;192mb\033[38;2;197;202;195mk\033[38;2;194;196;192mb\033[38;2;175;180;177mq\033[38;2;144;155;152mQ\033[38;2;109;128;123mX\033[38;2;71;101;94mr\033[38;2;46;89;78m?\033[38;2;39;91;78m?\033[38;2;43;100;89mf\033[38;2;47;108;99mj\033[38;2;51;115;104mr\033[38;2;54;117;105mx\033[38;2;52;115;104mr\033[38;2;54;117;106mx\033[38;2;56;118;103mx\033[38;2;56;119;101mx\033[38;2;58;121;102mx\033[38;2;58;123;104mn\033[38;2;58;124;105mnn\033[38;2;58;124;104mn\033[38;2;57;127;105mn\033[38;2;48;104;86mf\033[38;2;20;54;42m!\033[38;2;37;74;60m_\033[38;2;65;120;101mn\033[38;2;62;130;107mn\033[38;2;62;127;107mn\033[38;2;64;127;109mu\033[38;2;64;128;110muu\033[38;2;63;128;110mu\033[38;2;63;128;111mu\033[38;2;64;128;107mn\033[38;2;59;129;107mn\033[38;2;52;133;116mu\033[38;2;46;152;137mc\033[38;2;48;190;178mC\033[38;2;64;227;218mm\033[38;2;72;237;231mq\033[38;2;57;212;206mO\033[38;2;46;167;155mX\033[38;2;50;134;116mu\033[38;2;57;122;103mx\033[38;2;52;122;101mx\033[38;2;55;121;103mx\033[38;2;56;120;103mx\033[38;2;56;119;103mx\033[38;2;47;111;95mj\033[38;2;41;98;83m1\033[38;2;26;63;54mi\033[38;2;11;30;25m,\033[38;2;7;17;13m'\033[38;2;1;12;8m.\033[38;2;2;15;10m.\033[38;2;3;15;11m.\033[38;2;6;27;15m \033[38;2;46;132;94mr\033[38;2;58;219;159mL\033[38;2;44;214;151mJ\033[38;2;49;193;139mY\033[38;2;57;160;119mc\033[38;2;69;142;111mv\033[38;2;82;130;107mv\033[38;2;98;127;110mc\033[38;2;124;144;130mU\033[38;2;144;171;155m0\033[38;2;167;196;179mq\033[38;2;196;219;200ma\033[38;2;221;237;216mM\033[38;2;237;251;227m8\033[38;2;234;250;226m&\033[38;2;204;242;216m#\033[38;2;142;216;195mp\033[38;2;68;168;154mU\033[38;2;28;88;82m-\033[38;2;7;12;13m'\033[38;2;22;61;54mi\033[38;2;41;138;132mu\033[38;2;37;131;123mn\033[38;2;39;125;118mx\033[38;2;38;160;145mz\033[38;2;32;206;193mL\033[38;2;14;246;240mm\033[38;2;46;172;171mU\033[38;2;217;219;216m*\033[38;2;254;255;255m \033[38;2;255;255;254m \033[38;2;220;249;247m8\033[38;2;120;234;228mb\033[38;2;129;246;242ma\033[38;2;100;233;227md\033[38;2;126;228;219mb\033[38;2;208;240;229mM\033[38;2;254;255;253m \033[38;2;255;255;255m \033[38;2;255;254;255m  \033[38;2;255;255;254m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m           \033[38;2;232;234;233m&\033[38;2;167;174;169mm\033[38;2;78;104;93mx\033[38;2;37;86;74m-\033[38;2;41;99;88mf\033[38;2;71;119;108mn\033[38;2;107;144;134mU\033[38;2;144;167;158m0\033[38;2;173;186;178mq\033[38;2;197;202;196mk\033[38;2;184;188;184md\033[38;2;152;157;154m0\033[38;2;117;131;127mY\033[38;2;84;111;104mn\033[38;2;51;93;84mf\033[38;2;41;95;83m1\033[38;2;43;106;91mf\033[38;2;49;116;98mr\033[38;2;52;119;101mr\033[38;2;54;116;99mr\033[38;2;52;116;97mr\033[38;2;50;113;95mr\033[38;2;48;108;91mj\033[38;2;53;114;97mr\033[38;2;56;122;104mx\033[38;2;59;117;102mx\033[38;2;26;61;53mi\033[38;2;39;80;69m-\033[38;2;65;127;107mn\033[38;2;59;126;105mn\033[38;2;58;126;104mn\033[38;2;60;125;104mn\033[38;2;60;125;105mn\033[38;2;61;126;106mn\033[38;2;62;126;108mn\033[38;2;61;126;108mn\033[38;2;61;127;103mn\033[38;2;62;127;106mn\033[38;2;64;127;110mu\033[38;2;61;125;109mn\033[38;2;57;126;108mn\033[38;2;56;129;112mn\033[38;2;46;147;132mv\033[38;2;47;179;165mU\033[38;2;62;214;205mO\033[38;2;62;228;223mw\033[38;2;53;190;180mC\033[38;2;51;132;117mu\033[38;2;56;120;100mx\033[38;2;57;121;104mx\033[38;2;55;120;106mx\033[38;2;54;119;104mx\033[38;2;53;117;100mr\033[38;2;43;104;88mf\033[38;2;42;95;82m1\033[38;2;24;59;49mi\033[38;2;10;27;21m,\033[38;2;4;15;11m'\033[38;2;1;19;13m'\033[38;2;3;23;17m'\033[38;2;2;24;14m'\033[38;2;4;20;6m'\033[38;2;39;126;91mj\033[38;2;63;247;182mZ\033[38;2;55;246;179mO\033[38;2;46;187;140mY\033[38;2;44;141;111mn\033[38;2;44;132;106mx\033[38;2;40;114;95mj\033[38;2;42;100;88mf\033[38;2;37;92;83m?\033[38;2;35;83;75m-\033[38;2;38;82;75m-\033[38;2;46;87;80m?\033[38;2;66;105;99mr\033[38;2;93;137;128mX\033[38;2;110;168;149mC\033[38;2;114;178;160mQ\033[38;2;94;185;168mQ\033[38;2;68;196;182mQ\033[38;2;42;147;143mc\033[38;2;37;91;90m1\033[38;2;35;136;123mn\033[38;2;35;182;172mU\033[38;2;37;187;183mJ\033[38;2;39;152;143mc\033[38;2;33;192;177mJ\033[38;2;23;249;245mw\033[38;2;36;172;173mY\033[38;2;188;200;198mk\033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;171;242;237m*\033[38;2;149;247;245mo\033[38;2;187;243;242mM\033[38;2;210;246;244m&\033[38;2;252;254;253m \033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m             \033[38;2;246;246;243mB\033[38;2;176;184;180mq\033[38;2;84;107;102mn\033[38;2;42;83;73m-\033[38;2;33;79;66m_\033[38;2;45;81;70m-\033[38;2;70;91;84mj\033[38;2;103;115;108mv\033[38;2;122;125;120mX\033[38;2;144;143;137mC\033[38;2;176;173;168mw\033[38;2;196;191;187mb\033[38;2;183;182;178mp\033[38;2;154;159;155m0\033[38;2;104;120;113mc\033[38;2;70;97;87mj\033[38;2;55;82;74m?\033[38;2;63;82;79m1\033[38;2;73;89;84mj\033[38;2;88;99;95mx\033[38;2;109;117;114mc\033[38;2;126;142;137mJ\033[38;2;92;122;112mv\033[38;2;40;71;62m_\033[38;2;31;64;57m~\033[38;2;56;118;102mx\033[38;2;52;127;106mn\033[38;2;57;126;107mn\033[38;2;58;124;106mn\033[38;2;57;125;105mn\033[38;2;57;126;98mx\033[38;2;56;125;99mx\033[38;2;56;126;104mn\033[38;2;56;125;106mn\033[38;2;59;124;105mn\033[38;2;61;125;107mn\033[38;2;62;126;109mn\033[38;2;61;126;109mn\033[38;2;60;124;107mn\033[38;2;62;123;104mn\033[38;2;59;122;104mn\033[38;2;55;125;109mn\033[38;2;52;132;117mu\033[38;2;50;147;129mv\033[38;2;55;153;135mz\033[38;2;50;134;121mu\033[38;2;59;153;139mz\033[38;2;50;135;121mu\033[38;2;52;118;108mx\033[38;2;56;116;104mx\033[38;2;54;118;101mx\033[38;2;41;105;89mf\033[38;2;44;101;86mf\033[38;2;37;79;67m_\033[38;2;12;36;28m;\033[38;2;3;16;12m'\033[38;2;1;16;11m.\033[38;2;1;18;12m'\033[38;2;4;17;10m'\033[38;2;3;4;0m \033[38;2;31;115;79m1\033[38;2;65;249;179mZ\033[38;2;51;229;162mQ\033[38;2;51;175;133mX\033[38;2;39;122;99mr\033[38;2;55;136;117mu\033[38;2;53;134;116mu\033[38;2;52;128;114mn\033[38;2;51;123;111mn\033[38;2;48;117;106mr\033[38;2;46;109;99mj\033[38;2;42;98;88mf\033[38;2;35;85;76m-\033[38;2;27;73;67m+\033[38;2;24;65;63m~\033[38;2;29;69;68m+\033[38;2;40;96;88m1\033[38;2;43;121;112mx\033[38;2;35;167;164mX\033[38;2;47;183;173mJ\033[38;2;36;110;109mj\033[38;2;33;125;118mx\033[38;2;26;182;173mY\033[38;2;30;221;210m0\033[38;2;18;233;230mO\033[38;2;15;253;248mw\033[38;2;34;154;158mz\033[38;2;194;200;198mk\033[38;2;255;255;255m \033[38;2;251;253;253m \033[38;2;150;239;233ma\033[38;2;201;251;250m&\033[38;2;255;255;253m \033[38;2;255;255;255m \033[38;2;255;255;254m  \033[38;2;255;255;255m           ");
  $display("\033[38;2;255;255;255m               \033[38;2;248;247;246m@\033[38;2;199;199;196mk\033[38;2;191;191;189mb\033[38;2;225;224;222mM\033[38;2;245;244;244mB\033[38;2;255;254;254m \033[38;2;252;251;251m@\033[38;2;243;242;242mB\033[38;2;232;231;230mW\033[38;2;225;222;220m#\033[38;2;220;216;215m*\033[38;2;246;242;240mB\033[38;2;255;255;255m \033[38;2;242;240;239m8\033[38;2;234;232;231mW\033[38;2;243;241;240m8\033[38;2;251;249;249m@\033[38;2;255;255;255m   \033[38;2;248;247;247m@\033[38;2;217;216;216m*\033[38;2;176;187;184mp\033[38;2;113;142;132mU\033[38;2;70;114;99mx\033[38;2;54;107;91mj\033[38;2;54;115;99mr\033[38;2;57;121;105mx\033[38;2;58;124;105mn\033[38;2;60;126;107mn\033[38;2;61;125;108mn\033[38;2;61;124;108mn\033[38;2;60;124;107mnn\033[38;2;60;125;107mn\033[38;2;59;123;106mn\033[38;2;58;122;106mn\033[38;2;57;122;103mx\033[38;2;57;121;104mx\033[38;2;58;120;104mx\033[38;2;58;120;102mx\033[38;2;58;119;102mx\033[38;2;56;118;103mx\033[38;2;56;121;107mx\033[38;2;54;132;115mu\033[38;2;50;127;110mn\033[38;2;55;117;102mx\033[38;2;56;118;103mx\033[38;2;55;118;103mx\033[38;2;42;103;87mf\033[38;2;34;80;68m_\033[38;2;26;56;47mi\033[38;2;11;27;21m,\033[38;2;4;8;7m..\033[38;2;5;13;10m.\033[38;2;5;7;4m.\033[38;2;18;55;34ml\033[38;2;66;185;137mU\033[38;2;44;158;114mv\033[38;2;37;120;90mj\033[38;2;49;127;104mx\033[38;2;52;135;116mu\033[38;2;53;133;116mu\033[38;2;54;129;114mn\033[38;2;54;125;111mn\033[38;2;52;120;107mx\033[38;2;49;115;103mr\033[38;2;50;110;100mr\033[38;2;50;108;99mj\033[38;2;47;109;98mj\033[38;2;45;106;95mj\033[38;2;43;96;89mf\033[38;2;39;83;79m?\033[38;2;29;66;64m+\033[38;2;19;47;47ml\033[38;2;19;50;45m!\033[38;2;21;95;87m?\033[38;2;43;146;142mc\033[38;2;38;98;95mf\033[38;2;41;126;114mx\033[38;2;26;188;176mU\033[38;2;20;246;244mm\033[38;2;28;251;248mw\033[38;2;24;92;96m?\033[38;2;160;156;157mO\033[38;2;249;247;246m@\033[38;2;255;255;252m \033[38;2;149;237;235ma\033[38;2;212;250;250m&\033[38;2;255;253;254m \033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                                       \033[38;2;244;242;242mB\033[38;2;205;208;207ma\033[38;2;157;174;169mm\033[38;2;112;143;135mU\033[38;2;74;116;104mn\033[38;2;54;102;89mj\033[38;2;53;110;95mr\033[38;2;53;119;102mx\033[38;2;55;124;106mn\033[38;2;56;125;107mn\033[38;2;56;124;106mn\033[38;2;58;123;106mn\033[38;2;58;122;104mx\033[38;2;57;122;97mx\033[38;2;57;122;100mx\033[38;2;55;120;103mx\033[38;2;54;119;101mx\033[38;2;55;119;102mx\033[38;2;55;120;104mx\033[38;2;55;119;103mx\033[38;2;54;119;100mx\033[38;2;54;135;113mu\033[38;2;51;134;113mn\033[38;2;51;113;98mr\033[38;2;43;94;81m1\033[38;2;25;60;50mi\033[38;2;13;31;25m,\033[38;2;6;13;11m'\033[38;2;3;6;5m \033[38;2;1;6;4m \033[38;2;2;8;6m.\033[38;2;3;8;9m.\033[38;2;4;10;6m.\033[38;2;49;103;78mf\033[38;2;44;119;94mj\033[38;2;49;116;100mr\033[38;2;56;135;117mu\033[38;2;52;135;117mu\033[38;2;54;129;114mn\033[38;2;55;127;113mn\033[38;2;54;125;111mn\033[38;2;53;119;107mx\033[38;2;51;114;103mr\033[38;2;49;111;100mr\033[38;2;52;109;100mr\033[38;2;52;106;98mj\033[38;2;46;103;94mj\033[38;2;44;102;92mf\033[38;2;43;100;91mf\033[38;2;42;98;89mf\033[38;2;39;93;85m1\033[38;2;35;84;77m-\033[38;2;29;71;65m+\033[38;2;20;53;49m!\033[38;2;16;47;45ml\033[38;2;25;49;48m!\033[38;2;17;36;32m;\033[38;2;47;143;133mv\033[38;2;42;211;198mQ\033[38;2;27;124;120mr\033[38;2;11;35;33m;\033[38;2;27;97;86m?\033[38;2;85;188;184m0\033[38;2;140;226;222mk\033[38;2;100;234;231md\033[38;2;191;248;246mW\033[38;2;255;255;254m \033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m                         \033[38;2;255;255;254m \033[38;2;255;255;255m    \033[38;2;255;255;254m \033[38;2;252;252;249m@\033[38;2;249;249;246m@\033[38;2;244;244;242mB\033[38;2;240;239;239m8\033[38;2;221;218;218m#\033[38;2;150;149;148mQ\033[38;2;93;101;97mn\033[38;2;134;148;142mC\033[38;2;184;192;188md\033[38;2;219;221;220m#\033[38;2;241;239;239m8\033[38;2;244;241;241mB\033[38;2;227;228;224mM\033[38;2;210;210;207mo\033[38;2;170;182;175mw\033[38;2;123;151;139mJ\033[38;2;86;128;113mv\033[38;2;63;118;100mx\033[38;2;59;123;105mn\033[38;2;59;127;108mn\033[38;2;58;126;103mn\033[38;2;59;123;98mx\033[38;2;57;122;101mx\033[38;2;55;121;105mx\033[38;2;57;119;105mx\033[38;2;53;120;104mx\033[38;2;51;121;105mx\033[38;2;51;122;105mx\033[38;2;49;121;102mr\033[38;2;46;119;99mr\033[38;2;38;100;85m1\033[38;2;23;66;55m~\033[38;2;8;34;25m,\033[38;2;4;13;10m.\033[38;2;4;6;5m.\033[38;2;2;7;5m \033[38;2;4;5;3m \033[38;2;2;7;1m \033[38;2;0;8;4m \033[38;2;4;10;9m.\033[38;2;29;61;52mi\033[38;2;48;108;93mj\033[38;2;52;125;110mn\033[38;2;54;127;114mn\033[38;2;53;126;112mn\033[38;2;52;126;111mn\033[38;2;54;122;110mn\033[38;2;52;120;108mx\033[38;2;52;116;104mr\033[38;2;50;110;100mr\033[38;2;47;109;98mj\033[38;2;49;108;99mj\033[38;2;49;106;97mj\033[38;2;47;104;95mj\033[38;2;44;101;92mf\033[38;2;42;101;91mf\033[38;2;42;99;90mf\033[38;2;41;94;86m1\033[38;2;41;92;85m1\033[38;2;36;93;84m?\033[38;2;32;90;83m?\033[38;2;30;83;77m-\033[38;2;29;75;70m_\033[38;2;22;60;57mi\033[38;2;13;27;27m,\033[38;2;12;23;25m,\033[38;2;16;37;35mI\033[38;2;2;11;11m.\033[38;2;4;9;10m.\033[38;2;2;54;49ml\033[38;2;16;169;165mz\033[38;2;25;231;232mZ\033[38;2;21;237;237mZ\033[38;2;143;243;243mo\033[38;2;249;255;255m \033[38;2;255;254;255m \033[38;2;254;254;254m \033[38;2;253;255;255m \033[38;2;252;250;251m@\033[38;2;244;244;243mB\033[38;2;243;242;241mB\033[38;2;245;243;242mB\033[38;2;255;255;255m   \033[38;2;254;255;255m \033[38;2;255;255;255m   ");
  $display("\033[38;2;255;255;255m                         \033[38;2;254;255;252m \033[38;2;231;232;225mW\033[38;2;179;182;174mq\033[38;2;132;147;138mC\033[38;2;109;138;127mY\033[38;2;102;135;124mX\033[38;2;91;126;115mc\033[38;2;85;122;109mv\033[38;2;78;114;103mn\033[38;2;72;107;98mx\033[38;2;59;95;87mf\033[38;2;39;88;76m?\033[38;2;48;108;92mj\033[38;2;51;111;95mj\033[38;2;50;105;90mj\033[38;2;58;109;96mr\033[38;2;71;117;106mn\033[38;2;81;123;113mv\033[38;2;94;127;116mc\033[38;2;113;141;130mU\033[38;2;133;154;146mL\033[38;2;147;165;158m0\033[38;2;145;159;150mQ\033[38;2;106;125;116mz\033[38;2;55;87;76m1\033[38;2;40;84;70m-\033[38;2;50;101;84mf\033[38;2;53;113;97mr\033[38;2;54;120;103mx\033[38;2;57;121;103mx\033[38;2;57;122;106mn\033[38;2;51;125;105mx\033[38;2;50;121;102mx\033[38;2;46;108;91mj\033[38;2;35;87;72m-\033[38;2;21;59;49mi\033[38;2;9;31;27m,\033[38;2;2;15;12m.\033[38;2;2;9;7m.\033[38;2;2;8;6m.\033[38;2;0;6;4m \033[38;2;0;6;2m \033[38;2;4;27;21m \033[38;2;23;86;75m_\033[38;2;30;106;94mf\033[38;2;35;103;90mf\033[38;2;54;124;108mn\033[38;2;51;118;103mr\033[38;2;48;109;97mj\033[38;2;47;101;93mf\033[38;2;46;96;84m1\033[38;2;45;94;80m1\033[38;2;44;93;86m1\033[38;2;41;91;85m1\033[38;2;43;89;83m?\033[38;2;43;89;84m1\033[38;2;45;97;90mf\033[38;2;49;105;96mj\033[38;2;48;105;96mj\033[38;2;44;101;92mf\033[38;2;42;99;90mf\033[38;2;39;95;86m1\033[38;2;38;94;85m1\033[38;2;35;90;81m?\033[38;2;31;86;78m-\033[38;2;33;88;82m?\033[38;2;37;87;83m?\033[38;2;35;82;79m-\033[38;2;32;79;77m-\033[38;2;29;75;75m_\033[38;2;27;66;67m+\033[38;2;17;39;38mI\033[38;2;5;9;7m.\033[38;2;5;9;11m.\033[38;2;3;7;9m.\033[38;2;5;23;20m \033[38;2;4;91;85m_\033[38;2;18;200;195mJ\033[38;2;18;245;248mm\033[38;2;71;245;242md\033[38;2;201;254;253m&\033[38;2;253;254;255m \033[38;2;250;255;254m \033[38;2;146;202;198mp\033[38;2;54;116;111mx\033[38;2;38;60;59m~\033[38;2;37;40;42m!\033[38;2;38;36;37ml\033[38;2;100;98;99mn\033[38;2;245;244;245mB\033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;255;255;255m   ");
  $display("\033[38;2;255;255;255m                         \033[38;2;255;255;254m \033[38;2;253;253;252m \033[38;2;237;238;236m&\033[38;2;190;196;193mb\033[38;2;139;155;151mQ\033[38;2;84;118;109mu\033[38;2;47;93;83m1\033[38;2;37;94;83m?\033[38;2;40;106;93mf\033[38;2;46;114;102mr\033[38;2;52;116;105mx\033[38;2;53;118;106mx\033[38;2;53;119;104mx\033[38;2;56;120;105mx\033[38;2;54;120;106mx\033[38;2;52;118;105mxx\033[38;2;51;117;103mr\033[38;2;50;116;99mr\033[38;2;49;114;97mr\033[38;2;47;113;96mj\033[38;2;47;111;95mj\033[38;2;50;109;97mj\033[38;2;56;110;98mr\033[38;2;55;106;92mj\033[38;2;51;99;85mf\033[38;2;48;97;85mf\033[38;2;48;104;90mf\033[38;2;55;118;100mx\033[38;2;56;121;102mx\033[38;2;49;115;97mr\033[38;2;37;99;81m1\033[38;2;25;72;58m~\033[38;2;13;43;34mI\033[38;2;4;23;18m \033[38;2;0;15;10m.\033[38;2;1;15;9m.\033[38;2;3;12;9m.\033[38;2;2;6;6m \033[38;2;1;9;5m.\033[38;2;13;36;23m;\033[38;2;34;83;60m_\033[38;2;37;107;85mf\033[38;2;42;150;131mv\033[38;2;55;174;159mU\033[38;2;42;124;110mx\033[38;2;24;59;52mi\033[38;2;34;57;54m~\033[38;2;36;76;65m_\033[38;2;36;82;72m-\033[38;2;41;89;80m?\033[38;2;46;97;87mf\033[38;2;49;103;94mj\033[38;2;49;105;97mj\033[38;2;51;106;98mj\033[38;2;51;107;98mj\033[38;2;50;106;97mj\033[38;2;49;106;97mj\033[38;2;48;105;96mj\033[38;2;46;103;94mj\033[38;2;44;101;92mf\033[38;2;41;99;87m1\033[38;2;41;98;88m1\033[38;2;39;97;89m1\033[38;2;36;93;86m?\033[38;2;35;88;84m?\033[38;2;36;85;82m?\033[38;2;35;82;80m-\033[38;2;34;78;77m-\033[38;2;32;74;73m_\033[38;2;22;69;67m~\033[38;2;22;66;62m~\033[38;2;20;53;51m!\033[38;2;17;44;44ml\033[38;2;18;34;33m;\033[38;2;5;15;15m'\033[38;2;1;46;40mI\033[38;2;10;117;111mf\033[38;2;20;204;202mC\033[38;2;31;243;237mm\033[38;2;105;248;245mk\033[38;2;216;253;254m8\033[38;2;255;254;254m \033[38;2;217;238;237mW\033[38;2;73;143;138mz\033[38;2;0;64;59m!\033[38;2;0;34;36m,\033[38;2;15;31;32m;\033[38;2;0;2;4m \033[38;2;113;109;109mc\033[38;2;252;252;250m@\033[38;2;255;255;255m    ");
  $display("\033[38;2;255;255;255m                              \033[38;2;250;249;248m@\033[38;2;215;217;214m*\033[38;2;163;172;167mm\033[38;2;102;124;118mz\033[38;2;61;96;88mj\033[38;2;44;91;80m?\033[38;2;40;98;84m1\033[38;2;43;109;93mj\033[38;2;50;113;99mr\033[38;2;54;115;104mx\033[38;2;54;116;106mx\033[38;2;53;118;106mx\033[38;2;52;119;106mx\033[38;2;53;118;105mx\033[38;2;54;118;104mx\033[38;2;55;120;106mx\033[38;2;56;122;107mn\033[38;2;56;123;105mx\033[38;2;57;123;106mn\033[38;2;56;122;106mx\033[38;2;56;122;107mn\033[38;2;52;122;104mx\033[38;2;53;115;99mr\033[38;2;45;99;84mf\033[38;2;31;77;64m_\033[38;2;16;51;42ml\033[38;2;4;29;22m \033[38;2;1;16;9m.\033[38;2;2;15;9m.\033[38;2;2;16;10m.\033[38;2;3;14;8m.\033[38;2;1;14;5m.\033[38;2;8;33;20m,\033[38;2;25;83;61m+\033[38;2;49;142;106mn\033[38;2;53;144;106mu\033[38;2;38;108;79m1\033[38;2;38;103;82m1\033[38;2;51;122;103mx\033[38;2;45;99;85mf\033[38;2;13;32;25m,\033[38;2;21;42;37mI\033[38;2;44;105;96mj\033[38;2;42;133;122mn\033[38;2;42;136;129mu\033[38;2;42;129;121mn\033[38;2;46;118;109mx\033[38;2;50;110;100mr\033[38;2;49;107;97mj\033[38;2;49;106;97mj\033[38;2;48;105;96mj\033[38;2;47;104;95mj\033[38;2;47;101;93mf\033[38;2;44;99;90mf\033[38;2;43;97;89mff\033[38;2;42;96;89m1\033[38;2;39;93;88m1\033[38;2;38;91;87m1\033[38;2;36;89;86m?\033[38;2;37;88;85m?\033[38;2;35;85;82m?\033[38;2;33;82;79m-\033[38;2;32;79;76m-\033[38;2;28;77;74m_\033[38;2;21;67;64m~\033[38;2;18;63;58mi\033[38;2;18;66;60m~\033[38;2;15;60;57mi\033[38;2;34;76;74m_\033[38;2;29;60;56m~\033[38;2;3;20;18m'\033[38;2;6;61;54m!\033[38;2;8;130;123mr\033[38;2;22;210;208mL\033[38;2;40;246;243mq\033[38;2;165;251;250m#\033[38;2;219;251;248m8\033[38;2;244;255;253m@\033[38;2;250;252;251m@\033[38;2;151;203;199mp\033[38;2;17;77;75m+\033[38;2;5;23;24m \033[38;2;2;9;8m.\033[38;2;5;5;4m \033[38;2;168;165;161mZ\033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m        \033[38;2;254;255;254m \033[38;2;255;255;255m                         \033[38;2;233;232;231mW\033[38;2;185;188;187md\033[38;2;124;137;133mU\033[38;2;68;93;86mj\033[38;2;35;66;58m+\033[38;2;28;67;58m~\033[38;2;30;82;69m_\033[38;2;36;95;80m?\033[38;2;40;96;82m1\033[38;2;40;94;80m?\033[38;2;38;92;79m?\033[38;2;37;85;75m-\033[38;2;36;76;69m_\033[38;2;34;72;63m+\033[38;2;34;70;62m+\033[38;2;34;70;63m+\033[38;2;32;67;61m+\033[38;2;26;61;52mi\033[38;2;17;42;35mI\033[38;2;8;22;17m \033[38;2;3;11;7m.\033[38;2;3;9;7m.\033[38;2;3;10;7m.\033[38;2;1;11;7m.\033[38;2;1;12;7m.\033[38;2;5;22;15m'\033[38;2;17;66;45m!\033[38;2;35;134;94mr\033[38;2;59;196;143mU\033[38;2;58;188;137mY\033[38;2;32;121;86mf\033[38;2;31;96;77m?\033[38;2;48;117;103mr\033[38;2;57;126;110mn\033[38;2;43;86;75m?\033[38;2;12;27;23m,\033[38;2;29;60;53mi\033[38;2;53;113;100mr\033[38;2;37;138;123mn\033[38;2;41;183;174mU\033[38;2;67;225;219mm\033[38;2;47;194;184mC\033[38;2;36;140;131mu\033[38;2;41;111;100mj\033[38;2;42;103;92mf\033[38;2;43;101;92mf\033[38;2;43;100;91mf\033[38;2;40;97;88m1\033[38;2;39;93;85m1\033[38;2;40;93;85m1\033[38;2;41;94;86m1\033[38;2;42;95;87m1\033[38;2;40;92;84m1\033[38;2;39;91;84m?\033[38;2;38;90;85m?\033[38;2;37;90;85m?\033[38;2;35;90;85m?\033[38;2;33;86;82m?\033[38;2;31;82;79m-\033[38;2;30;81;78m-\033[38;2;28;78;77m_\033[38;2;28;72;71m_\033[38;2;24;64;62m~\033[38;2;21;57;57mi\033[38;2;20;61;60mi\033[38;2;16;58;57mi\033[38;2;45;105;100mj\033[38;2;24;56;57mi\033[38;2;5;27;23m \033[38;2;6;77;69m~\033[38;2;14;141;139mn\033[38;2;22;217;215mQ\033[38;2;48;250;247mp\033[38;2;68;248;246md\033[38;2;83;225;220mq\033[38;2;213;237;236mW\033[38;2;255;255;255m \033[38;2;140;151;147mL\033[38;2;4;11;6m.\033[38;2;2;4;9m.\033[38;2;1;1;1m \033[38;2;141;138;136mC\033[38;2;255;255;255m    ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;254;255;251m \033[38;2;236;245;235m \033[38;2;218;238;220m \033[38;2;215;242;218m \033[38;2;216;242;219m  \033[38;2;216;242;218m \033[38;2;216;242;219m    \033[38;2;216;242;220m \033[38;2;217;243;220m \033[38;2;216;242;220m  \033[38;2;216;243;219m \033[38;2;215;243;218m   \033[38;2;213;243;219m \033[38;2;217;241;218m \033[38;2;213;243;217m \033[38;2;223;241;227m \033[38;2;250;252;250m \033[38;2;255;255;255m     \033[38;2;247;246;246mB\033[38;2;207;205;205ma\033[38;2;142;144;144mL\033[38;2;71;83;80mf\033[38;2;24;44;39ml\033[38;2;8;32;25m,\033[38;2;9;39;28m;\033[38;2;12;42;31m;\033[38;2;10;32;27m,\033[38;2;6;17;17m'\033[38;2;0;4;7m \033[38;2;0;2;6m  \033[38;2;0;1;5m \033[38;2;0;2;3m \033[38;2;1;3;2m \033[38;2;2;3;0m \033[38;2;1;4;0m \033[38;2;1;9;3m \033[38;2;10;21;14m \033[38;2;15;59;41m!\033[38;2;34;121;88mj\033[38;2;49;185;134mX\033[38;2;58;221;162mQ\033[38;2;51;187;137mY\033[38;2;35;123;93mj\033[38;2;29;97;74m-\033[38;2;41;111;87mf\033[38;2;46;114;97mj\033[38;2;40;97;88m1\033[38;2;35;73;66m_\033[38;2;20;40;38mI\033[38;2;45;82;79m?\033[38;2;49;113;100mr\033[38;2;43;112;96mj\033[38;2;40;124;111mx\033[38;2;39;149;138mv\033[38;2;41;158;153mz\033[38;2;45;166;157mX\033[38;2;34;130;119mx\033[38;2;37;105;96mf\033[38;2;40;101;91mf\033[38;2;41;100;90mf\033[38;2;42;99;90mf\033[38;2;41;97;88m1\033[38;2;43;96;88m11\033[38;2;42;95;87m1\033[38;2;40;93;84m1\033[38;2;39;92;82m?\033[38;2;39;92;83m?\033[38;2;37;90;83m?\033[38;2;35;88;82m?\033[38;2;32;85;81m-\033[38;2;31;82;78m-\033[38;2;32;81;78m-\033[38;2;30;78;76m_\033[38;2;27;74;74m_\033[38;2;27;72;71m+\033[38;2;25;67;65m~\033[38;2;20;60;60mi\033[38;2;19;58;60mi\033[38;2;22;58;59mi\033[38;2;16;68;67m~\033[38;2;57;141;134mc\033[38;2;12;32;36m;\033[38;2;10;44;38mI\033[38;2;10;87;81m_\033[38;2;14;150;144mu\033[38;2;20;229;222mO\033[38;2;74;252;253mb\033[38;2;84;241;240md\033[38;2;65;190;186mQ\033[38;2;226;236;237m&\033[38;2;255;255;255m \033[38;2;143;139;136mC\033[38;2;2;5;6m \033[38;2;10;11;13m'\033[38;2;204;202;199mh\033[38;2;255;255;255m    ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;254;254m \033[38;2;255;254;255m \033[38;2;132;206;138mO\033[38;2;22;180;38mf\033[38;2;15;193;34mf\033[38;2;14;193;36mj\033[38;2;14;193;37mj\033[38;2;14;193;38mj\033[38;2;14;193;39mj\033[38;2;16;192;39mj\033[38;2;17;191;39mj\033[38;2;16;192;40mj\033[38;2;14;192;41mj\033[38;2;14;193;41mj\033[38;2;13;193;40mj\033[38;2;13;193;41mj\033[38;2;14;193;39mj\033[38;2;14;194;38mj\033[38;2;14;193;38mj\033[38;2;14;193;39mj\033[38;2;13;193;43mj\033[38;2;15;193;38mj\033[38;2;11;193;35mf\033[38;2;56;188;72mv\033[38;2;224;243;225m \033[38;2;255;255;255m  \033[38;2;255;254;255m  \033[38;2;255;255;255m    \033[38;2;254;252;253m \033[38;2;211;209;210mo\033[38;2;135;133;134mJ\033[38;2;59;62;60m_\033[38;2;11;15;13m'\033[38;2;0;0;0m \033[38;2;0;2;2m \033[38;2;2;6;8m.\033[38;2;1;6;7m \033[38;2;1;5;7m \033[38;2;0;3;5m \033[38;2;0;2;3m \033[38;2;2;2;4m \033[38;2;0;11;8m.\033[38;2;16;51;38ml\033[38;2;32;114;82mf\033[38;2;47;183;133mX\033[38;2;56;219;160mL\033[38;2;56;211;154mC\033[38;2;43;160;115mv\033[38;2;23;89;63m_\033[38;2;14;50;36mI\033[38;2;23;52;43m!\033[38;2;24;55;46m!\033[38;2;24;57;47m!\033[38;2;29;64;56m~\033[38;2;39;80;74m-\033[38;2;40;98;87m1\033[38;2;45;112;98mj\033[38;2;47;113;102mr\033[38;2;43;109;98mj\033[38;2;45;110;97mj\033[38;2;41;99;84m1\033[38;2;22;60;52mi\033[38;2;30;70;64m+\033[38;2;43;102;93mf\033[38;2;40;104;95mf\033[38;2;41;100;94mf\033[38;2;39;100;92mf\033[38;2;41;98;91mf\033[38;2;44;98;89mf\033[38;2;42;99;88mf\033[38;2;39;95;86m1\033[38;2;38;94;85m1\033[38;2;38;94;86m1\033[38;2;37;93;84m?\033[38;2;37;90;81m?\033[38;2;35;87;80m?\033[38;2;33;86;80m-\033[38;2;31;82;79m-\033[38;2;30;79;78m-\033[38;2;30;78;77m_\033[38;2;29;77;76m_\033[38;2;29;75;74m_\033[38;2;29;73;74m_\033[38;2;28;71;74m_\033[38;2;27;70;70m+\033[38;2;24;66;65m~\033[38;2;24;54;57mi\033[38;2;13;52;51m!\033[38;2;12;35;38m;\033[38;2;31;114;108mj\033[38;2;43;126;127mn\033[38;2;7;28;29m,\033[38;2;12;68;60mi\033[38;2;13;99;98m?\033[38;2;17;174;168mX\033[38;2;41;242;235mw\033[38;2;62;253;252md\033[38;2;32;217;217m0\033[38;2;93;142;139mY\033[38;2;248;249;244m@\033[38;2;255;252;254m \033[38;2;106;104;99mu\033[38;2;15;14;10m'\033[38;2;212;212;208mo\033[38;2;255;255;255m    ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;119;210;128m0\033[38;2;0;188;23m?\033[38;2;0;196;24m1\033[38;2;0;195;24m1\033[38;2;0;195;26m1\033[38;2;0;194;28m1\033[38;2;0;194;29m1\033[38;2;0;195;29m1\033[38;2;0;195;27m1\033[38;2;0;194;21m?\033[38;2;0;194;16m?\033[38;2;0;194;17m?\033[38;2;0;193;20m?\033[38;2;0;194;21m?\033[38;2;0;196;24m1\033[38;2;0;196;25m1\033[38;2;0;197;23m1\033[38;2;0;197;22m1\033[38;2;0;196;22m1\033[38;2;0;197;18m?\033[38;2;0;195;18m?\033[38;2;41;191;61mn\033[38;2;221;241;226m \033[38;2;255;255;255m           \033[38;2;254;252;254m \033[38;2;208;205;207ma\033[38;2;136;132;135mJ\033[38;2;59;57;57m_\033[38;2;15;15;15m  \033[38;2;24;24;24m;\033[38;2;35;36;36ml\033[38;2;48;48;52m~\033[38;2;59;59;61m_\033[38;2;74;87;80mf\033[38;2;96;130;113mc\033[38;2;101;163;136mJ\033[38;2;95;173;141mJ\033[38;2;91;152;126mX\033[38;2;54;82;68m?\033[38;2;15;17;15m \033[38;2;0;0;0m \033[38;2;0;2;1m \033[38;2;1;7;6m \033[38;2;9;22;17m \033[38;2;22;43;38ml\033[38;2;28;64;56m~\033[38;2;32;79;70m_\033[38;2;39;93;84m1\033[38;2;40;100;89mf\033[38;2;41;101;90mf\033[38;2;38;90;82m?\033[38;2;36;67;63m+\033[38;2;12;29;26m,\033[38;2;32;62;60m~\033[38;2;50;98;92mf\033[38;2;42;97;89mf\033[38;2;39;98;91mf\033[38;2;41;98;92mf\033[38;2;41;98;90mf\033[38;2;37;94;86m1\033[38;2;37;92;83m?\033[38;2;37;90;83m?\033[38;2;36;87;82m?\033[38;2;32;84;79m-\033[38;2;32;83;78m-\033[38;2;29;80;75m_\033[38;2;29;78;76m_\033[38;2;30;80;77m-\033[38;2;31;80;77m-\033[38;2;29;78;75m_\033[38;2;29;78;74m_\033[38;2;29;78;76m_\033[38;2;28;76;79m_\033[38;2;28;75;79m_\033[38;2;29;74;78m_\033[38;2;29;68;77m_\033[38;2;29;62;69m+\033[38;2;19;52;51m!\033[38;2;16;37;34mI\033[38;2;7;26;25m,\033[38;2;7;14;15m'\033[38;2;9;82;75m+\033[38;2;63;200;196m0\033[38;2;10;48;47ml\033[38;2;15;50;44ml\033[38;2;15;64;69m~\033[38;2;12;102;100m?\033[38;2;21;188;182mU\033[38;2;22;249;245mw\033[38;2;20;252;251mw\033[38;2;28;139;136mu\033[38;2;182;181;179mq\033[38;2;255;255;255m \033[38;2;204;199;191mk\033[38;2;127;122;113mX\033[38;2;254;254;252m \033[38;2;255;255;255m \033[38;2;255;255;254m \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;118;212;130m0\033[38;2;0;189;25m?\033[38;2;0;195;26m1\033[38;2;2;195;28m1\033[38;2;2;195;29m1\033[38;2;2;194;28m1\033[38;2;3;194;28m1\033[38;2;4;194;25m1\033[38;2;11;194;36mf\033[38;2;63;203;78mz\033[38;2;78;205;93mY\033[38;2;76;206;93mY\033[38;2;75;206;98mY\033[38;2;37;197;60mn\033[38;2;1;196;25m1\033[38;2;0;197;26m1\033[38;2;0;197;27m1\033[38;2;0;196;29m1\033[38;2;2;195;29m1\033[38;2;2;196;23m1\033[38;2;0;194;23m1\033[38;2;43;190;64mn\033[38;2;219;242;225m \033[38;2;255;255;255m \033[38;2;242;248;241m \033[38;2;219;239;220m \033[38;2;240;250;241m    \033[38;2;239;250;241m \033[38;2;240;250;241m   \033[38;2;240;251;243m \033[38;2;242;254;242m \033[38;2;240;247;236m \033[38;2;245;244;244m \033[38;2;227;225;225m \033[38;2;227;224;224m \033[38;2;238;236;236m \033[38;2;248;246;246m \033[38;2;255;254;253m \033[38;2;255;255;255m     \033[38;2;252;248;250m@\033[38;2;243;241;241m8\033[38;2;211;209;208mo\033[38;2;151;148;147mQ\033[38;2;83;86;84mj\033[38;2;34;38;37ml\033[38;2;3;9;7m.\033[38;2;0;0;0m \033[38;2;0;0;1m \033[38;2;1;10;8m.\033[38;2;9;23;18m \033[38;2;16;33;27m;\033[38;2;18;34;30m;\033[38;2;16;30;29m;\033[38;2;20;39;38mI\033[38;2;29;64;59m~\033[38;2;40;92;86m1\033[38;2;40;96;88m1\033[38;2;38;96;88m1\033[38;2;38;98;90m1\033[38;2;38;81;79m-\033[38;2;27;59;55mi\033[38;2;39;84;77m-\033[38;2;34;88;82m?\033[38;2;35;87;84m?\033[38;2;36;87;83m?\033[38;2;34;85;82m?\033[38;2;32;83;80m-\033[38;2;32;82;79m-\033[38;2;34;82;84m-\033[38;2;34;82;83m-\033[38;2;32;80;79m-\033[38;2;30;78;75m_\033[38;2;27;77;76m_\033[38;2;27;76;74m_\033[38;2;28;76;74m_\033[38;2;26;73;70m+\033[38;2;23;65;62m~\033[38;2;20;52;53m!\033[38;2;18;39;41mI\033[38;2;8;20;21m \033[38;2;6;11;13m'\033[38;2;4;7;10m.\033[38;2;1;20;19m'\033[38;2;25;153;145mv\033[38;2;45;221;213mO\033[38;2;11;48;51ml\033[38;2;15;33;35m;\033[38;2;13;47;49ml\033[38;2;16;60;60mi\033[38;2;10;111;103m1\033[38;2;26;217;212mQ\033[38;2;11;254;255mw\033[38;2;30;211;211mQ\033[38;2;101;134;130mX\033[38;2;253;253;250m \033[38;2;232;228;225mW\033[38;2;237;235;231m&\033[38;2;255;255;255m \033[38;2;255;255;254m  \033[38;2;255;255;255m  ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;116;212;129m0\033[38;2;0;190;24m?\033[38;2;0;196;26m1\033[38;2;0;196;28m1\033[38;2;0;196;27m1\033[38;2;1;197;26m1\033[38;2;1;196;25m1\033[38;2;4;192;24m1\033[38;2;40;188;65mn\033[38;2;212;238;212m#\033[38;2;255;255;255m  \033[38;2;255;254;255m \033[38;2;124;211;138mO\033[38;2;1;190;26m1\033[38;2;2;197;23m1\033[38;2;3;195;23m1\033[38;2;4;193;30m1\033[38;2;4;193;34mf\033[38;2;2;195;27m1\033[38;2;0;194;24m1\033[38;2;42;191;65mn\033[38;2;219;241;226m \033[38;2;255;255;255m \033[38;2;168;225;177m \033[38;2;24;188;42mj\033[38;2;34;199;57mn\033[38;2;36;199;59mn\033[38;2;35;198;58mn\033[38;2;36;199;60mn\033[38;2;35;197;58mnn\033[38;2;35;199;60mnn\033[38;2;36;197;60mn\033[38;2;35;198;55mn\033[38;2;55;180;66m \033[38;2;148;178;142m \033[38;2;172;182;169m \033[38;2;188;199;188mb\033[38;2;188;198;190mb\033[38;2;180;192;186md\033[38;2;181;192;188md\033[38;2;179;188;185mp\033[38;2;177;185;183mp\033[38;2;183;189;186md\033[38;2;176;177;173mw\033[38;2;196;191;189mb\033[38;2;242;238;236m8\033[38;2;255;255;255m    \033[38;2;239;239;239m8\033[38;2;195;195;195mk\033[38;2;132;132;132mU\033[38;2;74;73;73m1\033[38;2;33;31;31mI\033[38;2;10;9;7m.\033[38;2;0;0;0m \033[38;2;0;1;2m \033[38;2;5;13;14m'\033[38;2;11;26;25m,\033[38;2;19;43;41ml\033[38;2;25;55;53mi\033[38;2;32;71;69m_\033[38;2;37;83;79m-\033[38;2;31;63;59m~\033[38;2;16;37;33m;\033[38;2;35;72;66m_\033[38;2;40;91;83m?\033[38;2;34;90;83m?\033[38;2;33;88;82m?\033[38;2;35;85;82m?\033[38;2;34;84;81m-\033[38;2;33;83;80m-\033[38;2;32;83;79m-\033[38;2;33;82;82m-\033[38;2;33;80;79m-\033[38;2;32;76;74m_\033[38;2;31;73;72m_\033[38;2;25;70;70m+\033[38;2;24;64;64m~\033[38;2;25;57;59mi\033[38;2;18;42;44ml\033[38;2;11;27;30m,\033[38;2;6;17;19m'\033[38;2;4;8;11m.\033[38;2;3;5;7m.\033[38;2;2;5;7m \033[38;2;5;6;8m.\033[38;2;10;83;77m+\033[38;2;34;233;227mZ\033[38;2;33;190;186mJ\033[38;2;4;32;32m,\033[38;2;5;16;19m'\033[38;2;6;17;16m'\033[38;2;12;31;29m;\033[38;2;7;55;49ml\033[38;2;22;174;166mX\033[38;2;14;254;252mw\033[38;2;18;245;238mm\033[38;2;69;137;138mz\033[38;2;245;242;240mB\033[38;2;255;255;255m       ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;114;211;128mQ\033[38;2;0;189;23m?\033[38;2;1;195;26m1\033[38;2;2;195;27m1\033[38;2;0;195;28m1\033[38;2;0;196;29m1\033[38;2;4;194;28m1\033[38;2;3;194;25m1\033[38;2;37;190;63mn\033[38;2;208;239;210m#\033[38;2;255;255;255m \033[38;2;255;255;253m \033[38;2;255;253;255m \033[38;2;126;209;140mO\033[38;2;0;191;24m?\033[38;2;0;198;23m1\033[38;2;1;197;25m1\033[38;2;2;194;31m1\033[38;2;2;194;33mf\033[38;2;1;196;27m1\033[38;2;0;195;23m1\033[38;2;41;193;59mn\033[38;2;221;241;225m \033[38;2;252;254;251m \033[38;2;97;200;113mJ\033[38;2;0;192;19m?\033[38;2;0;196;24m1\033[38;2;0;194;23m1\033[38;2;0;195;22m1\033[38;2;0;194;22m1\033[38;2;7;196;35mf\033[38;2;2;195;28m1\033[38;2;0;194;20m?\033[38;2;0;195;23m1\033[38;2;0;192;29m1\033[38;2;0;196;20m1\033[38;2;3;191;28m1\033[38;2;145;213;155m \033[38;2;178;186;178mq\033[38;2;77;114;98mn\033[38;2;37;91;75m?\033[38;2;36;87;75m-\033[38;2;32;88;75m-\033[38;2;30;88;77m-\033[38;2;34;88;78m-\033[38;2;27;59;52mi\033[38;2;106;110;105mv\033[38;2;213;210;210mo\033[38;2;249;247;247m@\033[38;2;255;254;254m \033[38;2;255;255;253m \033[38;2;255;255;252m \033[38;2;255;255;254m \033[38;2;255;255;255m  \033[38;2;250;247;247m@\033[38;2;198;196;196mk\033[38;2;172;169;168mm\033[38;2;148;144;144mL\033[38;2;99;96;97mn\033[38;2;44;43;44mi\033[38;2;3;3;3m \033[38;2;1;0;0m \033[38;2;2;1;2m \033[38;2;3;5;6m \033[38;2;9;12;13m'\033[38;2;7;18;15m'\033[38;2;6;8;9m.\033[38;2;25;54;48m!\033[38;2;33;87;78m-\033[38;2;35;88;81m?\033[38;2;34;88;79m?\033[38;2;32;87;79m-\033[38;2;30;84;78m-\033[38;2;32;82;78m-\033[38;2;33;74;74m_\033[38;2;29;65;66m+\033[38;2;28;61;61m~\033[38;2;23;52;52m!\033[38;2;21;45;46ml\033[38;2;19;39;40mI\033[38;2;11;26;28m,\033[38;2;8;21;22m \033[38;2;6;14;14m'\033[38;2;3;8;9m.\033[38;2;2;5;8m.\033[38;2;0;5;6m \033[38;2;0;5;5m \033[38;2;2;6;5m \033[38;2;2;8;6m.\033[38;2;6;51;45ml\033[38;2;29;195;186mJ\033[38;2;28;251;249mq\033[38;2;21;104;107mf\033[38;2;6;13;13m'\033[38;2;4;8;12m.\033[38;2;3;7;6m.\033[38;2;6;29;27m,\033[38;2;17;114;109mf\033[38;2;27;228;223mO\033[38;2;9;255;255mw\033[38;2;24;205;203mL\033[38;2;126;159;158mQ\033[38;2;251;251;249m@\033[38;2;254;254;255m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;112;211;127mQ\033[38;2;0;189;23m?\033[38;2;3;195;25m1\033[38;2;3;194;26m1\033[38;2;0;196;29m1\033[38;2;1;195;31m1\033[38;2;4;193;30m1\033[38;2;0;195;22m1\033[38;2;42;186;60mn\033[38;2;204;239;209m*\033[38;2;255;253;253m \033[38;2;253;254;253m \033[38;2;253;254;251m \033[38;2;123;210;137m0\033[38;2;1;188;27m1\033[38;2;1;198;25m1\033[38;2;0;197;28m1\033[38;2;3;194;29m1\033[38;2;3;194;27m1\033[38;2;1;197;25m1\033[38;2;0;195;25m1\033[38;2;43;191;60mn\033[38;2;224;243;227m \033[38;2;221;244;222m \033[38;2;33;190;55mx\033[38;2;0;196;24m1\033[38;2;1;196;30m1\033[38;2;1;196;25m1\033[38;2;0;199;26m1\033[38;2;4;190;27m1\033[38;2;120;214;131m0\033[38;2;72;203;89mX\033[38;2;0;193;21m?\033[38;2;3;196;23m1\033[38;2;3;194;30m1\033[38;2;2;194;25m1\033[38;2;0;194;21m?\033[38;2;81;197;100m \033[38;2;251;255;252m \033[38;2;239;240;241m8\033[38;2;189;198;196mb\033[38;2;170;180;176mw\033[38;2;156;165;162mO\033[38;2;149;158;158m0\033[38;2;135;148;144mC\033[38;2;148;148;147mQ\033[38;2;255;251;255m \033[38;2;255;255;255m      \033[38;2;255;255;253m \033[38;2;254;255;254m \033[38;2;251;248;251m@\033[38;2;222;213;217m@\033[38;2;162;150;155m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;255;255;255m@\033[38;2;1;2;2m \033[38;2;2;5;7m \033[38;2;7;12;12m'\033[38;2;9;23;20m \033[38;2;15;33;30m;\033[38;2;19;39;35mI\033[38;2;19;42;37mI\033[38;2;16;39;33mI\033[38;2;13;32;28m;\033[38;2;11;23;23m,\033[38;2;11;18;21m \033[38;2;8;13;16m'\033[38;2;5;9;12m.\033[38;2;3;6;9m.\033[38;2;2;5;8m.\033[38;2;0;4;7m \033[38;2;0;4;5m \033[38;2;0;5;4m \033[38;2;1;6;4m \033[38;2;1;8;6m.\033[38;2;3;9;6m.\033[38;2;1;9;6m.\033[38;2;1;12;6m.\033[38;2;4;50;36mI\033[38;2;32;174;165mX\033[38;2;19;255;251mw\033[38;2;32;200;198mL\033[38;2;8;36;37m;\033[38;2;5;15;7m.\033[38;2;0;13;8m.\033[38;2;4;43;37m;\033[38;2;20;148;141mu\033[38;2;23;240;238mm\033[38;2;7;255;255mw\033[38;2;22;221;218m0\033[38;2;68;121;121mu\033[38;2;235;232;233m&\033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;112;211;126mQ\033[38;2;0;190;24m?\033[38;2;2;195;25m1\033[38;2;2;196;26m1\033[38;2;0;198;27m1\033[38;2;1;196;27m1\033[38;2;3;195;26m1\033[38;2;3;196;21m1\033[38;2;13;193;32mf\033[38;2;51;202;70mv\033[38;2;67;201;78mz\033[38;2;67;200;84mz\033[38;2;63;201;82mz\033[38;2;30;197;50mx\033[38;2;3;195;23m1\033[38;2;1;196;21m1\033[38;2;1;196;27m1\033[38;2;4;193;32mf\033[38;2;3;194;29m1\033[38;2;2;198;23m1\033[38;2;0;196;18m?\033[38;2;46;187;66mn\033[38;2;232;244;234m \033[38;2;155;221;159m \033[38;2;4;191;23m1\033[38;2;1;196;26m1\033[38;2;1;195;32mf\033[38;2;1;195;26m1\033[38;2;0;195;26m1\033[38;2;29;187;46mr\033[38;2;213;241;215m \033[38;2;159;220;163m \033[38;2;6;187;35mf\033[38;2;2;196;28m1\033[38;2;3;195;27m1\033[38;2;3;196;22m1\033[38;2;0;195;27m1\033[38;2;23;188;48mr\033[38;2;201;237;207m \033[38;2;255;255;255m   \033[38;2;247;255;250m \033[38;2;166;232;175m \033[38;2;116;221;132m0\033[38;2;113;221;126m0\033[38;2;107;216;122mQ\033[38;2;105;212;116mL\033[38;2;105;211;120mL\033[38;2;102;212;122mL\033[38;2;103;212;117mL\033[38;2;99;214;107mC\033[38;2;116;210;135m0\033[38;2;233;246;236m8\033[38;2;255;255;255m \033[38;2;209;241;211m \033[38;2;9;193;29mm\033[38;2;9;193;29m0\033[38;2;9;193;29mL\033[38;2;9;193;29mj\033[38;2;9;193;29m!\033[38;2;9;193;29mi\033[38;2;9;193;29mi\033[38;2;9;193;29mi\033[38;2;9;193;29m+\033[38;2;9;193;29m!\033[38;2;255;255;255m@\033[38;2;2;1;6m \033[38;2;1;1;3m \033[38;2;1;0;0m \033[38;2;1;1;0m  \033[38;2;1;0;0m \033[38;2;1;1;0m \033[38;2;1;1;1m \033[38;2;0;1;2m \033[38;2;1;2;4m \033[38;2;2;1;6m \033[38;2;1;2;7m \033[38;2;0;4;7m  \033[38;2;3;5;9m.\033[38;2;3;8;9m.\033[38;2;2;9;7m.\033[38;2;2;10;7m.\033[38;2;2;13;8m.\033[38;2;2;15;11m.\033[38;2;0;28;20m \033[38;2;10;76;61m~\033[38;2;36;187;173mU\033[38;2;28;251;254mq\033[38;2;26;232;229mZ\033[38;2;16;90;79m_\033[38;2;6;28;22m \033[38;2;0;40;29m,\033[38;2;13;104;93m?\033[38;2;26;202;197mC\033[38;2;12;255;252mw\033[38;2;11;255;255mw\033[38;2;19;213;205mL\033[38;2;64;119;118mu\033[38;2;211;211;207mo\033[38;2;255;255;255m \033[38;2;253;255;255m \033[38;2;255;255;254m \033[38;2;255;255;255m      ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;112;211;126mQ\033[38;2;0;190;24m?\033[38;2;3;195;26m1\033[38;2;3;194;28m1\033[38;2;0;197;26m1\033[38;2;0;197;23m1\033[38;2;1;196;24m1\033[38;2;2;195;30m1\033[38;2;1;193;32m1\033[38;2;0;193;22m?\033[38;2;0;195;15m?\033[38;2;0;195;17m?\033[38;2;0;195;20m?\033[38;2;0;194;20m?\033[38;2;1;193;23m1\033[38;2;0;195;24m1\033[38;2;0;197;25m1\033[38;2;0;196;27m1\033[38;2;0;196;24m1\033[38;2;0;190;26m1\033[38;2;15;183;36mf\033[38;2;139;210;146mZ\033[38;2;244;252;246m \033[38;2;81;197;90mX\033[38;2;0;194;23m1\033[38;2;5;193;29m1\033[38;2;0;196;31m1\033[38;2;7;193;23m1\033[38;2;0;193;22m?\033[38;2;88;197;107mU\033[38;2;255;254;255m \033[38;2;225;242;226m \033[38;2;41;188;62mn\033[38;2;1;196;24m1\033[38;2;2;197;25m1\033[38;2;2;196;25m1\033[38;2;1;195;26m1\033[38;2;1;188;25m?\033[38;2;136;214;147m \033[38;2;255;255;255m \033[38;2;255;254;253m \033[38;2;255;255;255m \033[38;2;159;226;170m \033[38;2;0;187;21m?\033[38;2;0;193;23m1\033[38;2;0;193;14m?\033[38;2;9;192;31mf\033[38;2;55;203;75mc\033[38;2;62;201;80mz\033[38;2;62;201;75mc\033[38;2;60;202;79mc\033[38;2;59;202;73mc\033[38;2;71;197;94mX\033[38;2;230;242;228m&\033[38;2;247;253;249m \033[38;2;61;198;80mc\033[38;2;0;189;19m?\033[38;2;0;193;19m?\033[38;2;0;194;22m1\033[38;2;39;206;59mu\033[38;2;70;212;88mX\033[38;2;68;212;94mY\033[38;2;72;211;92mY\033[38;2;51;188;66mu\033[38;2;9;193;29m?\033[38;2;9;193;29mi\033[38;2;255;255;255m@\033[38;2;2;3;4m \033[38;2;2;2;2m \033[38;2;1;2;4m \033[38;2;2;2;2m   \033[38;2;1;4;6m \033[38;2;0;4;6m \033[38;2;0;3;5m \033[38;2;0;4;7m \033[38;2;0;4;8m \033[38;2;1;5;8m \033[38;2;1;5;6m \033[38;2;2;5;5m \033[38;2;5;5;8m.\033[38;2;4;10;10m.\033[38;2;5;14;11m'\033[38;2;10;22;17m \033[38;2;13;31;26m,\033[38;2;19;46;37ml\033[38;2;31;80;66m_\033[38;2;37;127;107mr\033[38;2;33;141;130mu\033[38;2;32;140;131mu\033[38;2;25;93;82m-\033[38;2;4;18;10m'\033[38;2;8;43;37mI\033[38;2;36;172;162mX\033[38;2;20;254;247mw\033[38;2;7;255;255mw\033[38;2;13;255;253mw\033[38;2;22;176;175mY\033[38;2;75;112;112mn\033[38;2;218;217;214m*\033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;112;211;127mQ\033[38;2;0;190;24m?\033[38;2;3;195;27m1\033[38;2;1;195;29m1\033[38;2;0;196;28m1\033[38;2;2;195;27m1\033[38;2;4;195;25m1\033[38;2;2;196;24m1\033[38;2;4;194;29m1\033[38;2;18;194;39mj\033[38;2;24;194;44mr\033[38;2;22;195;43mr\033[38;2;23;194;43mr\033[38;2;28;190;48mr\033[38;2;28;190;50mr\033[38;2;23;195;45mr\033[38;2;22;197;43mr\033[38;2;27;194;50mr\033[38;2;46;194;67mu\033[38;2;94;203;108mJ\033[38;2;180;227;187mk\033[38;2;251;253;251m \033[38;2;207;236;211m \033[38;2;22;188;50mr\033[38;2;1;195;24m1\033[38;2;4;194;27m1\033[38;2;3;197;26m1\033[38;2;3;195;28m1\033[38;2;3;193;24m1\033[38;2;43;199;65mu\033[38;2;86;206;105mU\033[38;2;82;204;101mU\033[38;2;25;194;40mr\033[38;2;2;194;28m1\033[38;2;1;198;31mf\033[38;2;0;196;27m1\033[38;2;2;194;25m1\033[38;2;0;192;20m?\033[38;2;69;193;86mz\033[38;2;240;251;241m \033[38;2;255;254;255m \033[38;2;255;255;255m \033[38;2;146;221;156m \033[38;2;0;189;16m?\033[38;2;0;196;26m1\033[38;2;0;195;18m?\033[38;2;50;195;69mu\033[38;2;188;235;195ma\033[38;2;197;237;201mo\033[38;2;196;237;204mo\033[38;2;195;238;200mo\033[38;2;199;237;205mo\033[38;2;231;246;233m&\033[38;2;255;253;255m \033[38;2;239;251;243m \033[38;2;43;195;66mu\033[38;2;0;195;20m?\033[38;2;1;195;26m1\033[38;2;2;191;25m1\033[38;2;119;218;133m0\033[38;2;198;237;206mo\033[38;2;195;238;201mo\033[38;2;197;238;203mo\033[38;2;182;220;186mk\033[38;2;122;145;123mU\033[38;2;52;56;50m~\033[38;2;2;0;2m \033[38;2;0;0;0m       \033[38;2;0;1;0m \033[38;2;0;4;3m \033[38;2;2;5;4m \033[38;2;0;0;2m \033[38;2;1;0;0m  \033[38;2;1;1;0m \033[38;2;4;8;6m.\033[38;2;8;21;15m'\033[38;2;13;41;27m;\033[38;2;25;70;49m~\033[38;2;30;99;71m-\033[38;2;35;129;96mr\033[38;2;44;159;118mv\033[38;2;44;179;128mz\033[38;2;48;199;142mU\033[38;2;63;221;160mQ\033[38;2;44;147;99mn\033[38;2;42;119;84mj\033[38;2;22;66;49mi\033[38;2;16;66;62m~\033[38;2;27;179;174mY\033[38;2;29;225;224mO\033[38;2;27;138;138mu\033[38;2;114;132;125mX\033[38;2;240;236;233m&\033[38;2;255;255;255m           ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;114;213;127mQ\033[38;2;0;190;24m?\033[38;2;2;195;25m1\033[38;2;3;194;27m1\033[38;2;2;195;27m1\033[38;2;2;196;28m1\033[38;2;3;196;29mf\033[38;2;0;198;26m1\033[38;2;35;190;59mx\033[38;2;187;233;190mh\033[38;2;226;246;229m \033[38;2;226;246;226m  \033[38;2;226;245;227m  \033[38;2;226;246;227m  \033[38;2;227;246;228m \033[38;2;237;248;239m \033[38;2;255;255;255m   \033[38;2;135;215;148mm\033[38;2;1;190;28m1\033[38;2;4;194;29m1\033[38;2;2;196;31mf\033[38;2;5;194;26m1\033[38;2;0;197;28m1\033[38;2;0;193;22m?\033[38;2;0;191;16m?\033[38;2;0;192;13m?\033[38;2;0;191;13m?\033[38;2;0;193;14m?\033[38;2;0;195;25m1\033[38;2;3;195;25m1\033[38;2;2;195;25m1\033[38;2;1;196;26m1\033[38;2;0;197;24m1\033[38;2;20;186;44mj\033[38;2;193;231;199ma\033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;208;238;213m \033[38;2;57;195;77mv\033[38;2;9;193;29mf\033[38;2;7;194;27mf\033[38;2;6;192;32mf\033[38;2;8;190;33mf\033[38;2;8;192;31mf\033[38;2;8;191;32mf\033[38;2;5;193;27m1\033[38;2;4;194;31mf\033[38;2;41;194;63mn\033[38;2;206;239;213m#\033[38;2;252;254;253m \033[38;2;133;215;146mZ\033[38;2;24;192;41mj\033[38;2;6;193;32mf\033[38;2;5;194;31mf\033[38;2;7;192;34mf\033[38;2;8;191;36mf\033[38;2;8;191;32mf\033[38;2;4;194;30mf\033[38;2;8;193;30mf\033[38;2;20;201;42mr\033[38;2;109;199;115mC\033[38;2;164;165;168mZ\033[38;2;107;105;105mv\033[38;2;86;84;87mj\033[38;2;72;71;70m?\033[38;2;62;59;60m_\033[38;2;55;52;52m+\033[38;2;46;43;44mi\033[38;2;37;35;34ml\033[38;2;32;32;30mI\033[38;2;12;13;11m'\033[38;2;0;1;0m \033[38;2;17;40;29m;\033[38;2;25;70;49m~\033[38;2;38;102;74m?\033[38;2;47;136;99mx\033[38;2;53;165;121mc\033[38;2;58;181;134mY\033[38;2;56;194;142mU\033[38;2;59;207;151mC\033[38;2;59;219;158mL\033[38;2;55;225;164mQ\033[38;2;53;235;174m0\033[38;2;56;255;193mm\033[38;2;52;255;192mm\033[38;2;63;255;190mm\033[38;2;35;146;94mx\033[38;2;54;199;143mU\033[38;2;71;238;180mZ\033[38;2;37;103;74m?\033[38;2;0;8;2m \033[38;2;64;88;82mf\033[38;2;179;185;184mp\033[38;2;255;254;254m \033[38;2;255;255;255m \033[38;2;254;255;255m \033[38;2;255;255;255m          ");
  $display("\033[38;2;255;255;255m       \033[38;2;255;255;254m \033[38;2;255;255;255m \033[38;2;113;213;129mQ\033[38;2;0;189;24m?\033[38;2;1;196;28m1\033[38;2;1;196;30m1\033[38;2;2;195;30m1\033[38;2;1;194;28m1\033[38;2;0;195;25m1\033[38;2;0;190;23m?\033[38;2;80;193;99mY\033[38;2;241;250;240mB\033[38;2;255;255;255m         \033[38;2;252;255;255m \033[38;2;255;253;255m \033[38;2;241;249;240m \033[38;2;65;194;86mz\033[38;2;0;194;27m1\033[38;2;4;196;23m1\033[38;2;2;196;27m1\033[38;2;5;193;30mf\033[38;2;0;195;16m?\033[38;2;52;198;78mv\033[38;2;135;219;150mm\033[38;2;138;220;145mm\033[38;2;137;222;144mm\033[38;2;126;218;144mZ\033[38;2;29;192;52mx\033[38;2;0;194;22m1\033[38;2;4;195;27m1\033[38;2;2;195;29m1\033[38;2;0;196;28m1\033[38;2;1;188;27m1\033[38;2;124;209;132m0\033[38;2;255;255;254m \033[38;2;255;253;255m \033[38;2;255;255;255m \033[38;2;248;251;247m \033[38;2;211;241;219m \033[38;2;210;239;210m \033[38;2;204;241;210m \033[38;2;206;240;211m \033[38;2;208;241;208m \033[38;2;95;209;114mC\033[38;2;0;191;23m?\033[38;2;0;196;26m1\033[38;2;0;190;15m?\033[38;2;161;226;169md\033[38;2;255;255;255m \033[38;2;255;254;255m \033[38;2;230;245;231m \033[38;2;208;240;212m \033[38;2;208;241;211m \033[38;2;207;241;210m \033[38;2;209;241;211m \033[38;2;183;234;186mh\033[38;2;24;194;49mr\033[38;2;1;195;21m1\033[38;2;0;193;23m1\033[38;2;47;194;69mu\033[38;2;248;255;249m@\033[38;2;255;255;255m   \033[38;2;255;254;253m \033[38;2;252;252;250m@\033[38;2;248;248;246m@\033[38;2;243;242;240m8\033[38;2;240;240;238m8\033[38;2;206;207;205ma\033[38;2;120;124;120mX\033[38;2;61;94;78mf\033[38;2;27;85;61m_\033[38;2;25;80;59m+\033[38;2;22;71;53m~\033[38;2;17;60;45m!\033[38;2;12;52;39ml\033[38;2;10;46;34mI\033[38;2;9;44;32m;\033[38;2;8;48;33mI\033[38;2;8;54;36mI\033[38;2;6;67;42m!\033[38;2;43;159;117mv\033[38;2;60;255;191mm\033[38;2;59;232;169m0\033[38;2;26;156;108mn\033[38;2;63;204;170mL\033[38;2;33;145;113mn\033[38;2;58;114;87mr\033[38;2;132;137;126mU\033[38;2;239;235;233m&\033[38;2;255;255;255m              ");
  $display("\033[38;2;255;255;255m       \033[38;2;254;255;255m \033[38;2;254;255;253m \033[38;2;112;208;127mQ\033[38;2;0;186;14m-\033[38;2;0;191;20m?\033[38;2;0;193;17m?\033[38;2;0;193;18m?\033[38;2;3;190;24m1\033[38;2;20;189;39mj\033[38;2;84;203;103mU\033[38;2;209;239;219m#\033[38;2;255;254;255m \033[38;2;254;255;253m \033[38;2;254;255;255m       \033[38;2;255;254;254m \033[38;2;251;255;249m \033[38;2;255;253;255m \033[38;2;182;232;185mk\033[38;2;12;184;31m1\033[38;2;0;192;19m?\033[38;2;0;193;19m?\033[38;2;0;193;20m?\033[38;2;0;192;19m?\033[38;2;22;187;40mj\033[38;2;180;229;192mh\033[38;2;255;255;255m    \033[38;2;124;211;139mO\033[38;2;5;186;24m?\033[38;2;0;193;17m?\033[38;2;0;192;24m1\033[38;2;0;195;19m?\033[38;2;0;193;15m?\033[38;2;48;191;66mu\033[38;2;232;245;233m&\033[38;2;255;255;255m \033[38;2;193;231;198m \033[38;2;81;202;96mY\033[38;2;83;213;97mU\033[38;2;85;211;103mJ\033[38;2;85;211;102mU\033[38;2;88;209;100mU\033[38;2;85;212;100mU\033[38;2;36;198;58mn\033[38;2;0;193;23m1\033[38;2;0;193;16m?\033[38;2;4;188;29m1\033[38;2;187;231;191mh\033[38;2;252;255;254m \033[38;2;126;207;135m0\033[38;2;81;208;94mY\033[38;2;86;210;105mJ\033[38;2;85;211;103mJJ\033[38;2;86;211;104mJ\033[38;2;75;208;94mY\033[38;2;6;193;29mf\033[38;2;0;193;17m?\033[38;2;0;190;15m?\033[38;2;67;199;86mz\033[38;2;247;251;246m@\033[38;2;252;255;254m \033[38;2;254;254;252m \033[38;2;254;255;255m \033[38;2;255;255;255m       \033[38;2;222;218;218m#\033[38;2;123;117;118mX\033[38;2;23;20;20m,\033[38;2;0;0;0m \033[38;2;1;6;9m.\033[38;2;2;12;9m.\033[38;2;1;16;10m.\033[38;2;2;18;13m'\033[38;2;3;23;15m'\033[38;2;0;37;25m,\033[38;2;8;79;64m~\033[38;2;28;136;111mx\033[38;2;45;184;145mY\033[38;2;32;201;171mJ\033[38;2;30;174;163mX\033[38;2;46;131;122mn\033[38;2;113;135;130mY\033[38;2;218;216;214m*\033[38;2;255;255;255m                ");
  $display("\033[38;2;255;255;255m       \033[38;2;254;255;255m \033[38;2;254;252;253m \033[38;2;189;230;196ma\033[38;2;137;217;150mm\033[38;2;135;220;150mm\033[38;2;137;219;149mm\033[38;2;139;222;150mm\033[38;2;163;225;173md\033[38;2;208;239;213m#\033[38;2;249;252;249m@\033[38;2;255;254;255m  \033[38;2;254;255;254m \033[38;2;255;255;255m       \033[38;2;254;255;255m \033[38;2;255;254;254m \033[38;2;255;255;255m \033[38;2;177;224;178mb\033[38;2;89;205;103mU\033[38;2;88;211;105mJ\033[38;2;87;211;105mJ\033[38;2;90;211;106mJ\033[38;2;126;215;138mO\033[38;2;201;237;205m*\033[38;2;255;254;255m \033[38;2;253;254;255m \033[38;2;253;255;254m \033[38;2;253;254;254m \033[38;2;255;255;254m \033[38;2;245;252;245m \033[38;2;174;227;181mb\033[38;2;109;210;118mL\033[38;2;92;209;104mJ\033[38;2;89;210;100mJ\033[38;2;85;210;105mJ\033[38;2;101;201;125mC\033[38;2;217;238;218mM\033[38;2;254;254;255m \033[38;2;195;234;198m \033[38;2;70;203;90mX\033[38;2;69;207;84mX\033[38;2;68;208;85mX\033[38;2;69;208;85mX\033[38;2;69;207;85mX\033[38;2;69;207;87mX\033[38;2;75;208;92mY\033[38;2;79;208;95mY\033[38;2;89;208;104mJ\033[38;2;160;225;173md\033[38;2;250;252;248m \033[38;2;250;253;251m \033[38;2;123;210;138mO\033[38;2;63;207;82mz\033[38;2;70;206;88mX\033[38;2;68;207;86mX\033[38;2;68;208;86mXX\033[38;2;70;208;87mX\033[38;2;78;209;93mY\033[38;2;75;211;94mY\033[38;2;116;213;128m0\033[38;2;211;241;215m#\033[38;2;255;253;253m \033[38;2;253;255;254m \033[38;2;254;255;253m \033[38;2;254;255;255m \033[38;2;255;255;255m         \033[38;2;219;219;218m*\033[38;2;99;96;95mn\033[38;2;7;8;6m.\033[38;2;0;4;2m \033[38;2;2;15;13m'\033[38;2;1;19;11m'\033[38;2;1;46;32m;\033[38;2;17;124;112mj\033[38;2;41;196;187mC\033[38;2;34;183;181mU\033[38;2;29;142;134mu\033[38;2;51;124;117mn\033[38;2;121;145;146mJ\033[38;2;216;215;211m*\033[38;2;255;255;255m  \033[38;2;254;255;255m \033[38;2;255;255;255m               ");
  $display("\033[38;2;255;255;255m        \033[38;2;255;254;254m \033[38;2;255;255;255m        \033[38;2;254;255;254m \033[38;2;255;255;255m         \033[38;2;254;255;255m \033[38;2;255;255;255m            \033[38;2;255;254;255m \033[38;2;255;255;253m \033[38;2;255;255;255m        \033[38;2;253;255;255m \033[38;2;255;255;255m           \033[38;2;254;255;254m \033[38;2;255;254;255m \033[38;2;255;255;255m           \033[38;2;255;255;254m \033[38;2;254;255;255m  \033[38;2;255;255;255m        \033[38;2;255;255;254m \033[38;2;255;255;255m   \033[38;2;184;184;182mp\033[38;2;50;50;49m~\033[38;2;2;5;6m \033[38;2;13;68;60mi\033[38;2;37;148;140mv\033[38;2;36;156;153mz\033[38;2;30;110;109mj\033[38;2;70;105;101mx\033[38;2;147;155;151mQ\033[38;2;228;225;222mM\033[38;2;255;255;255m  \033[38;2;254;255;255m \033[38;2;255;255;255m                 ");
  $display("\033[38;2;255;255;255m                                                                                           \033[38;2;227;229;226mM\033[38;2;93;95;91mx\033[38;2;13;35;33m;\033[38;2;54;89;87mf\033[38;2;117;124;120mX\033[38;2;194;189;186md\033[38;2;245;244;242mB\033[38;2;255;255;255m                      ");
  $display("\033[38;2;255;255;255m                                                                                          \033[38;2;249;249;248m@\033[38;2;182;184;180mp\033[38;2;157;161;156mO\033[38;2;189;186;185md\033[38;2;236;232;231m&\033[38;2;255;255;255m                         ");
  $display("\033[38;2;255;255;255m                                                                                          \033[38;2;255;255;254m \033[38;2;255;255;255m                             ");
  $display("");
  $display ("--------------------------------------------------");
  $display("                  Congratulations!               ");
  $display("              execution cycles = %7d", total_latency);
  $display("              clock period = %4fns", CYCLE_clk1);
  $display ("--------------------------------------------------");
  $finish;	
endtask

task fail_task;
  $display("\033[0m                                                \033[38;2;255;255;255m$$$\033[38;2;247;247;247mB\033[38;2;241;241;241m%%\033[38;2;252;252;252m$\033[38;2;255;255;255m$$$\033[0m                                          \033[0m");
  $display("\033[0m                                             \033[38;2;255;255;255m$$\033[38;2;226;226;228mW\033[38;2;162;163;170mZ\033[38;2;116;119;128mz\033[38;2;98;102;113mu\033[38;2;95;99;112mn\033[38;2;94;98;111mn\033[38;2;93;96;107mx\033[38;2;95;99;106mn\033[38;2;122;125;127mX\033[38;2;167;167;169mm\033[38;2;231;231;229m&\033[38;2;255;255;255m$\033[0m                                        \033[0m");
  $display("\033[0m                                            \033[38;2;255;255;255m$\033[38;2;223;229;229mW\033[38;2;132;138;145mJ\033[38;2;60;66;81m?\033[38;2;72;77;91mt\033[38;2;107;112;123mc\033[38;2;145;148;157mQ\033[38;2;173;175;181mq\033[38;2;188;190;196mb\033[38;2;186;187;193md\033[38;2;123;126;137mY\033[38;2;30;36;53ml\033[38;2;30;35;52ml\033[38;2;67;71;85m1\033[38;2;159;158;161mO\033[38;2;251;251;248m@\033[38;2;255;255;255m$\033[0m                                      \033[0m");
  $display("\033[0m                                          \033[38;2;255;0;0mf\033[38;2;255;59;59mX\033[38;2;234;163;162md\033[38;2;110;60;68mt\033[38;2;80;57;69m?\033[38;2;189;197;202mk\033[38;2;249;255;253m$\033[38;2;255;255;255m$$$$$$\033[38;2;186;187;192md\033[38;2;37;43;58mi\033[38;2;30;36;54ml\033[38;2;27;30;45mI\033[38;2;189;186;184md\033[38;2;255;255;255m$\033[0m                                      \033[0m");
  $display("\033[0m                                \033[38;2;255;0;0mfffffff\033[38;2;255;1;1mf\033[38;2;255;2;2mj\033[38;2;255;0;0mff\033[38;2;255;69;69mU\033[38;2;254;65;65mY\033[38;2;249;51;52mz\033[38;2;255;34;33mu\033[38;2;244;84;86mJ\033[38;2;126;111;134mX\033[38;2;100;118;147mz\033[38;2;107;123;150mY\033[38;2;104;119;147mX\033[38;2;106;120;146mX\033[38;2;95;109;130mv\033[38;2;90;100;112mn\033[38;2;111;114;121mc\033[38;2;39;45;57mi\033[38;2;33;39;56m!\033[38;2;28;33;50ml\033[38;2;122;126;131mY\033[38;2;179;187;188mp\033[38;2;192;195;195mk\033[38;2;224;224;224mM\033[38;2;255;255;252m$\033[38;2;255;255;255m$\033[0m                                  \033[0m");
  $display("\033[0m                     \033[38;2;255;0;0mffff\033[0m    \033[38;2;255;0;0mfff\033[38;2;255;11;11mr\033[38;2;255;38;38mv\033[38;2;255;79;79mJ\033[38;2;255;109;109m0\033[38;2;255;141;141mq\033[38;2;255;173;173mh\033[38;2;255;195;195m*\033[38;2;255;210;210mW\033[38;2;255;215;215mW\033[38;2;255;154;154md\033[38;2;255;57;57mX\033[38;2;255;235;235m%%\033[38;2;255;255;255m$$\033[38;2;255;180;180ma\033[38;2;255;0;0mf\033[38;2;169;29;46mf\033[38;2;46;80;121mf\033[38;2;52;75;111mt\033[38;2;50;74;108mt\033[38;2;50;73;106m1\033[38;2;47;71;104m1\033[38;2;40;62;91m-\033[38;2;28;45;69mi\033[38;2;28;38;58m!\033[38;2;30;36;53ml\033[38;2;32;39;57m!\033[38;2;30;42;60m!\033[38;2;32;47;63mi\033[38;2;44;60;77m_\033[38;2;68;83;100mf\033[38;2;105;115;128mc\033[38;2;154;160;162mO\033[38;2;211;211;211mo\033[38;2;255;255;255m$$\033[0m                               \033[0m");
  $display("\033[0m           \033[38;2;255;0;0mffffff\033[0m   \033[38;2;255;0;0mff\033[38;2;255;21;21mn\033[38;2;255;14;14mr\033[38;2;255;2;2mj\033[38;2;255;0;0mff\033[0m  \033[38;2;255;0;0mff\033[38;2;255;143;143mp\033[38;2;255;225;225m8\033[38;2;255;252;252m$\033[38;2;255;255;255m$$$$\033[38;2;255;248;248m@\033[38;2;255;223;223m&\033[38;2;255;189;188mo\033[38;2;255;138;138mq\033[38;2;255;100;100mQ\033[38;2;255;251;251m$\033[38;2;255;255;255m$$\033[38;2;255;154;154md\033[38;2;255;0;0mf\033[38;2;127;49;72mf\033[38;2;48;81;119mf\033[38;2;54;80;115mf\033[38;2;50;79;113mt\033[38;2;51;75;108mt\033[38;2;53;73;107mt\033[38;2;54;74;109mt\033[38;2;52;74;109mt\033[38;2;47;67;101m?\033[38;2;35;49;71m~\033[38;2;27;36;51ml\033[38;2;27;36;50ml\033[38;2;28;36;52ml\033[38;2;26;35;53ml\033[38;2;25;34;53ml\033[38;2;25;34;54ml\033[38;2;29;44;62mi\033[38;2;56;72;87m?\033[38;2;116;127;136mY\033[38;2;190;192;194mb\033[38;2;255;255;255m$$\033[0m                             \033[0m");
  $display("\033[0m       \033[38;2;255;0;0mffff\033[38;2;255;15;15mx\033[38;2;255;45;45mc\033[38;2;255;77;77mJ\033[38;2;255;101;101mQ\033[38;2;255;79;79mJ\033[38;2;255;22;22mn\033[38;2;255;0;0mffff\033[38;2;255;110;110mO\033[38;2;255;233;233m%%\033[38;2;255;224;224m8\033[38;2;255;202;202m#\033[38;2;255;43;43mc\033[38;2;255;0;0mff\033[0m \033[38;2;255;0;0mff\033[38;2;255;70;70mU\033[38;2;255;210;210mWW\033[38;2;255;158;158mb\033[38;2;255;236;236m%%\033[38;2;255;255;255m$$\033[38;2;255;79;79mJ\033[38;2;248;9;10mj\033[38;2;225;9;15mf\033[38;2;255;0;0mf\033[38;2;255;131;131mw\033[38;2;255;255;255m$$\033[38;2;255;254;254m$\033[38;2;255;67;67mY\033[38;2;240;1;3mf\033[38;2;74;76;109mj\033[38;2;53;81;118mf\033[38;2;51;77;111mt\033[38;2;52;77;110mt\033[38;2;55;78;111mf\033[38;2;56;79;111mf\033[38;2;55;79;111mf\033[38;2;54;78;111mf\033[38;2;53;77;112mt\033[38;2;54;76;111mt\033[38;2;44;62;88m-\033[38;2;29;42;58m!\033[38;2;27;36;52ml\033[38;2;29;37;53ml\033[38;2;28;36;54ml\033[38;2;28;36;53ml\033[38;2;27;33;51ml\033[38;2;24;34;51ml\033[38;2;27;42;61m!\033[38;2;46;61;80m_\033[38;2;114;121;129mz\033[38;2;202;201;202mh\033[38;2;255;255;255m$$\033[0m                           \033[0m");
  $display("\033[0m    \033[38;2;255;0;0mfff\033[38;2;255;8;8mr\033[38;2;255;51;51mz\033[38;2;255;113;113mO\033[38;2;255;178;178ma\033[38;2;255;228;228m8\033[38;2;255;255;255m$$$$\033[38;2;255;222;222m&\033[38;2;255;58;58mX\033[38;2;255;4;4mj\033[38;2;255;84;84mC\033[38;2;255;153;153md\033[38;2;255;253;253m$\033[38;2;255;255;255m$$$\033[38;2;255;186;186mo\033[38;2;255;3;3mj\033[38;2;255;0;0mf\033[0m  \033[38;2;255;0;0mf\033[38;2;255;37;37mv\033[38;2;252;48;47mc\033[38;2;250;6;7mj\033[38;2;255;12;12mr\033[38;2;255;233;233m%%\033[38;2;255;255;255m$\033[38;2;255;246;246m@\033[38;2;255;31;30mu\033[38;2;208;14;23mf\033[38;2;169;37;54mj\033[38;2;255;2;2mj\033[38;2;255;203;203m#\033[38;2;255;255;255m$$\033[38;2;255;226;226m8\033[38;2;255;10;9mr\033[38;2;186;25;37mf\033[38;2;38;83;118mt\033[38;2;46;78;111mt\033[38;2;54;77;110mt\033[38;2;58;77;111mf\033[38;2;53;80;114mf\033[38;2;47;81;118mff\033[38;2;51;78;112mt\033[38;2;54;77;111mt\033[38;2;53;76;113mt\033[38;2;53;75;111mt\033[38;2;48;70;100m1\033[38;2;31;45;68mi\033[38;2;26;33;49ml\033[38;2;25;35;52ml\033[38;2;27;33;52ml\033[38;2;28;31;50ml\033[38;2;28;31;51ml\033[38;2;27;31;50ml\033[38;2;28;38;55ml\033[38;2;33;50;66mi\033[38;2;53;70;85m?\033[38;2;142;146;149mL\033[38;2;234;234;232m&\033[38;2;255;255;255m$\033[0m                          \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mff\033[38;2;255;22;22mn\033[38;2;255;75;75mJ\033[38;2;255;149;149mp\033[38;2;255;214;214mW\033[38;2;255;253;253m$\033[38;2;255;255;255m$$\033[38;2;255;236;236m%%\033[38;2;255;191;191m*\033[38;2;255;143;143mp\033[38;2;255;100;100mQ\033[38;2;255;68;68mY\033[38;2;255;46;46mc\033[38;2;255;7;7mj\033[38;2;255;115;115mO\033[38;2;255;255;255m$$$\033[38;2;255;249;249m@\033[38;2;255;255;255m$$$\033[38;2;255;117;117mZ\033[38;2;255;0;0mfff\033[38;2;255;214;214mW\033[38;2;202;218;222m*\033[38;2;119;115;134mX\033[38;2;231;1;5mt\033[38;2;255;53;53mz\033[38;2;255;254;254m$\033[38;2;255;255;255m$\033[38;2;255;220;220m&\033[38;2;255;6;5mj\033[38;2;184;29;43mf\033[38;2;214;13;21mf\033[38;2;255;37;36mv\033[38;2;255;247;247m@\033[38;2;255;255;255m$$\033[38;2;255;156;156mb\033[38;2;255;0;0mf\033[38;2;193;11;21m1\033[38;2;161;25;40m1\033[38;2;192;20;31mf\033[38;2;213;19;27mj\033[38;2;216;19;26mj\033[38;2;196;17;28mt\033[38;2;166;24;42mt\033[38;2;134;42;67mf\033[38;2;71;69;104mf\033[38;2;49;77;114mt\033[38;2;52;74;109mt\033[38;2;51;74;108mtt\033[38;2;50;72;105m1\033[38;2;34;47;70m~\033[38;2;27;32;51ml\033[38;2;26;35;53ml\033[38;2;25;36;52ml\033[38;2;27;34;52ml\033[38;2;26;32;50ml\033[38;2;26;30;49mI\033[38;2;25;32;48mI\033[38;2;33;50;64mi\033[38;2;36;57;73m+\033[38;2;84;95;106mx\033[38;2;202;204;203ma\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mf\033[38;2;255;6;6mj\033[38;2;255;195;195m*\033[38;2;255;255;255m$$$$\033[38;2;255;212;212mW\033[38;2;255;71;71mU\033[38;2;255;18;18mx\033[38;2;255;0;0mfffff\033[38;2;255;21;21mn\033[38;2;255;232;232m%%\033[38;2;255;255;255m$$\033[38;2;255;238;238mB\033[38;2;255;62;62mY\033[38;2;255;130;130mw\033[38;2;255;253;253m$\033[38;2;255;255;255m$\033[38;2;255;247;247m@\033[38;2;255;121;121mZ\033[38;2;255;103;103m0\033[38;2;255;65;65mY\033[38;2;255;35;35mv\033[38;2;187;38;49mr\033[38;2;116;55;81mf\033[38;2;255;0;0mf\033[38;2;255;137;137mq\033[38;2;255;255;255m$$\033[38;2;255;181;181ma\033[38;2;255;0;0mf\033[38;2;179;29;44mf\033[38;2;234;1;5mt\033[38;2;255;78;78mJ\033[38;2;255;255;255m$$$\033[38;2;255;121;121mZ\033[38;2;255;47;47mc\033[38;2;255;105;104m0\033[38;2;255;147;145mp\033[38;2;255;179;178ma\033[38;2;255;206;205mM\033[38;2;255;211;210mW\033[38;2;255;180;179ma\033[38;2;255;149;148mp\033[38;2;255;35;33mu\033[38;2;215;14;22mf\033[38;2;67;68;101mt\033[38;2;45;71;104m1\033[38;2;53;75;110mt\033[38;2;52;75;108mt\033[38;2;51;75;107mt\033[38;2;50;71;103m1\033[38;2;34;46;70m~\033[38;2;25;34;51ml\033[38;2;25;37;54ml\033[38;2;25;35;52mll\033[38;2;25;33;50ml\033[38;2;25;32;49mI\033[38;2;23;30;48mI\033[38;2;35;46;63mi\033[38;2;38;59;76m+\033[38;2;55;73;87m?\033[38;2;177;182;184mp\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mff\033[38;2;255;43;43mc\033[38;2;255;141;141mq\033[38;2;255;233;233m%%\033[38;2;255;255;255m$$\033[38;2;255;127;127mm\033[38;2;255;0;0mf\033[38;2;255;5;5mj\033[38;2;255;33;33mu\033[38;2;255;58;58mX\033[38;2;255;26;26mn\033[38;2;255;1;1mf\033[38;2;255;0;0mf\033[38;2;255;106;106m0\033[38;2;255;255;255m$$$\033[38;2;255;139;139mq\033[38;2;255;58;58mX\033[38;2;255;114;114mO\033[38;2;255;245;245m@\033[38;2;255;255;255m$$$$\033[38;2;255;188;188mo\033[38;2;255;15;14mr\033[38;2;229;1;6mt\033[38;2;206;11;20mt\033[38;2;255;6;5mj\033[38;2;255;219;219m&\033[38;2;255;255;255m$$\033[38;2;255;137;137mq\033[38;2;255;51;51mz\033[38;2;246;22;23mx\033[38;2;253;1;1mf\033[38;2;255;54;54mz\033[38;2;255;254;254m$\033[38;2;255;255;255m$$\033[38;2;255;248;248m@\033[38;2;255;254;254m$\033[38;2;255;255;255m$$$$\033[38;2;255;245;245m@\033[38;2;255;242;242mB\033[38;2;255;223;223m&\033[38;2;255;90;89mL\033[38;2;255;0;0mf\033[38;2;112;46;69m1\033[38;2;43;75;109m1\033[38;2;54;77;111mt\033[38;2;53;76;110mt\033[38;2;52;75;108mt\033[38;2;51;74;108mt\033[38;2;49;70;103m1\033[38;2;28;41;62m!\033[38;2;26;33;51ml\033[38;2;26;34;53ml\033[38;2;26;35;52mll\033[38;2;26;34;51ml\033[38;2;26;32;51ml\033[38;2;25;28;43mI\033[38;2;35;45;62mi\033[38;2;39;62;80m_\033[38;2;46;64;81m-\033[38;2;171;176;178mw\033[38;2;255;255;255m$\033[0m                       \033[0m");
  $display("\033[0m \033[38;2;255;0;0mff\033[38;2;255;1;1mf\033[38;2;255;37;37mv\033[38;2;255;54;54mz\033[38;2;255;219;219m&\033[38;2;255;255;255m$$\033[38;2;255;190;190mo\033[38;2;255;178;178ma\033[38;2;255;222;222m&\033[38;2;255;251;251m$\033[38;2;255;255;255m$\033[38;2;255;213;213mW\033[38;2;255;19;19mx\033[38;2;255;10;10mr\033[38;2;255;218;218m&\033[38;2;255;255;255m$$\033[38;2;255;250;250m@\033[38;2;255;252;252m$\033[38;2;255;255;255m$$$\033[38;2;255;240;240mB\033[38;2;255;255;255m$$\033[38;2;255;238;238mB\033[38;2;255;35;35mv\033[38;2;255;17;17mx\033[38;2;254;53;54mz\033[38;2;255;95;94mL\033[38;2;255;162;162mb\033[38;2;255;255;255m$$$$$\033[38;2;255;227;226m8\033[38;2;255;52;52mz\033[38;2;255;0;0mf\033[38;2;255;96;95mL\033[38;2;255;229;229m8\033[38;2;255;255;255m$$\033[38;2;255;240;239mB\033[38;2;255;195;194m*\033[38;2;255;130;129mw\033[38;2;255;83;83mC\033[38;2;251;49;49mc\033[38;2;237;32;33mn\033[38;2;234;30;33mn\033[38;2;223;20;25mj\033[38;2;192;20;31mf\033[38;2;120;46;68mt\033[38;2;81;82;95mj\033[38;2;54;75;105mt\033[38;2;54;76;112mt\033[38;2;53;77;112mt\033[38;2;53;75;110mt\033[38;2;52;74;106mt\033[38;2;53;75;108mt\033[38;2;44;63;88m-\033[38;2;24;36;53ml\033[38;2;27;37;53ml\033[38;2;26;35;52ml\033[38;2;25;34;51ml\033[38;2;26;35;52ml\033[38;2;25;34;51ml\033[38;2;25;32;49mI\033[38;2;25;30;46mI\033[38;2;36;49;66m~\033[38;2;40;63;80m_\033[38;2;44;63;78m_\033[38;2;171;175;177mw\033[38;2;255;255;255m$\033[0m                      \033[0m");
  $display("\033[0m \033[38;2;255;0;0mff\033[38;2;255;89;89mL\033[38;2;255;255;255m$$$$$$$\033[38;2;255;227;227m8\033[38;2;255;187;187mo\033[38;2;255;135;135mw\033[38;2;255;66;66mY\033[38;2;255;0;0mf\033[38;2;255;99;99mQ\033[38;2;255;255;255m$$\033[38;2;255;247;247m@\033[38;2;255;84;84mC\033[38;2;255;141;141mq\033[38;2;255;161;161mb\033[38;2;255;118;118mZ\033[38;2;255;77;77mJ\033[38;2;255;132;132mw\033[38;2;255;255;255m$$$\033[38;2;255;70;70mU\033[38;2;255;110;110mO\033[38;2;255;255;255m$$$\033[38;2;255;239;239mB\033[38;2;255;207;206mM\033[38;2;255;184;183mo\033[38;2;255;146;145mp\033[38;2;255;104;103m0\033[38;2;255;67;67mY\033[38;2;242;12;15mj\033[38;2;171;34;50mf\033[38;2;204;12;21mt\033[38;2;246;29;30mn\033[38;2;254;60;61mX\033[38;2;253;56;57mX\033[38;2;243;32;35mn\033[38;2;217;15;22mf\033[38;2;169;22;36m1\033[38;2;103;22;37m+\033[38;2;71;28;45mi\033[38;2;66;61;88m?\033[38;2;65;70;101mt\033[38;2;55;70;106mt\033[38;2;43;72;104m1\033[38;2;102;106;104mu\033[38;2;162;139;110mJ\033[38;2;61;77;97mt\033[38;2;53;73;103m1\033[38;2;55;73;102m1\033[38;2;52;76;111mt\033[38;2;52;75;108mt\033[38;2;49;72;104m1\033[38;2;47;68;101m1\033[38;2;34;46;69mi\033[38;2;26;36;52ml\033[38;2;27;37;54ml\033[38;2;24;31;49mI\033[38;2;25;33;51ml\033[38;2;25;34;51ml\033[38;2;25;35;52ml\033[38;2;26;32;50ml\033[38;2;25;32;47mI\033[38;2;37;54;69m~\033[38;2;39;61;77m_\033[38;2;45;64;80m-\033[38;2;200;202;202mh\033[38;2;255;255;255m$\033[0m                     \033[0m");
  $display("\033[0m \033[38;2;255;0;0mff\033[38;2;255;28;28mn\033[38;2;255;158;158mb\033[38;2;255;245;245m@\033[38;2;255;255;255m$$\033[38;2;255;189;189mo\033[38;2;255;90;90mL\033[38;2;255;43;43mc\033[38;2;255;13;13mr\033[38;2;255;0;0mfff\033[38;2;255;2;2mj\033[38;2;255;198;198m#\033[38;2;255;255;255m$$\033[38;2;255;204;204mM\033[38;2;255;0;0mfff\033[38;2;255;16;14mx\033[38;2;255;13;12mr\033[38;2;255;139;138mq\033[38;2;255;235;235m%%\033[38;2;255;224;223m8\033[38;2;255;124;122mm\033[38;2;255;4;4mj\033[38;2;255;8;8mr\033[38;2;255;112;111mO\033[38;2;255;126;125mm\033[38;2;255;74;73mU\033[38;2;246;33;35mu\033[38;2;218;19;26mj\033[38;2;193;21;33mf\033[38;2;185;20;34mt\033[38;2;138;38;59mt\033[38;2;111;52;79mt\033[38;2;83;70;103mf\033[38;2;49;82;121mf\033[38;2;49;70;107m1\033[38;2;74;57;88m1\033[38;2;92;52;79m1\033[38;2;91;58;85mt\033[38;2;76;65;98mt\033[38;2;57;76;111mf\033[38;2;34;61;87m_\033[38;2;22;41;61m!\033[38;2;45;69;97m?\033[38;2;50;77;113mt\033[38;2;44;71;109m1\033[38;2;61;75;97mt\033[38;2;133;123;102mz\033[38;2;207;181;139mw\033[38;2;220;193;156mb\033[38;2;88;89;98mr\033[38;2;55;74;94m1\033[38;2;115;108;101mv\033[38;2;51;71;98m1\033[38;2;52;74;107mt\033[38;2;53;73;104m1\033[38;2;37;54;83m+\033[38;2;40;56;82m_\033[38;2;27;35;52ml\033[38;2;25;37;54ml\033[38;2;25;33;49mI\033[38;2;23;32;47mI\033[38;2;26;34;52ml\033[38;2;26;34;51ml\033[38;2;26;33;51ml\033[38;2;25;30;47mI\033[38;2;26;36;52ml\033[38;2;37;60;74m+\033[38;2;34;55;76m+\033[38;2;80;92;102mr\033[38;2;237;237;234m8\033[38;2;255;255;255m$\033[0m                    \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mfff\033[38;2;255;219;219m&\033[38;2;255;255;255m$$\033[38;2;255;69;69mU\033[38;2;255;0;0mfff\033[0m  \033[38;2;255;0;0mf\033[38;2;255;1;1mf\033[38;2;255;89;89mL\033[38;2;255;206;206mM\033[38;2;255;208;208mM\033[38;2;255;84;84mC\033[38;2;253;0;0mf\033[38;2;255;85;85mC\033[38;2;255;255;255m$\033[38;2;168;164;176mm\033[38;2;162;40;57mj\033[38;2;217;13;20mf\033[38;2;239;31;34mn\033[38;2;235;25;29mx\033[38;2;199;17;28mf\033[38;2;121;57;84mj\033[38;2;107;61;91mj\033[38;2;156;29;46mt\033[38;2;154;32;51mt\033[38;2;119;49;75mf\033[38;2;80;68;103mf\033[38;2;57;80;119mf\033[38;2;49;84;125mj\033[38;2;49;85;125mj\033[38;2;48;85;122mf\033[38;2;52;83;122mf\033[38;2;54;81;120mf\033[38;2;55;77;114mf\033[38;2;47;70;106m1\033[38;2;40;65;94m-\033[38;2;47;77;108mt\033[38;2;50;80;114mf\033[38;2;50;79;114mf\033[38;2;48;72;102m1\033[38;2;29;39;63m!\033[38;2;46;62;90m-\033[38;2;49;73;108m1\033[38;2;52;67;100m1\033[38;2;103;99;101mn\033[38;2;189;165;131mO\033[38;2;233;212;169ma\033[38;2;246;226;187m#\033[38;2;250;230;191mM\033[38;2;181;169;153mm\033[38;2;50;63;90m-\033[38;2;143;126;112mY\033[38;2;121;115;115mz\033[38;2;49;67;96m?\033[38;2;57;75;106mt\033[38;2;40;55;81m+\033[38;2;34;48;70m~\033[38;2;28;39;60m!\033[38;2;25;36;53ml\033[38;2;26;34;52ml\033[38;2;23;30;49mI\033[38;2;26;34;52ml\033[38;2;26;34;51ml\033[38;2;26;34;52ml\033[38;2;26;33;49ml\033[38;2;23;30;46mI\033[38;2;30;45;60mi\033[38;2;38;60;76m+\033[38;2;32;53;73m~\033[38;2;129;136;142mJ\033[38;2;255;255;255m$\033[0m                    \033[0m");
  $display("\033[0m   \033[38;2;255;0;0mf\033[38;2;255;1;1mf\033[38;2;255;113;113mO\033[38;2;255;227;227m8\033[38;2;255;237;237mB\033[38;2;255;63;63mY\033[38;2;255;0;0mff\033[0m    \033[38;2;255;0;0mff\033[38;2;255;4;4mj\033[38;2;255;2;2mj\033[38;2;255;0;0mf\033[38;2;255;163;160mb\033[38;2;216;225;229mM\033[38;2;117;132;156mJ\033[38;2;51;77;116mf\033[38;2;52;88;126mj\033[38;2;61;83;121mj\033[38;2;78;77;112mj\033[38;2;74;78;114mj\033[38;2;57;86;127mr\033[38;2;52;87;128mj\033[38;2;48;81;120mf\033[38;2;47;84;120mf\033[38;2;48;86;126mj\033[38;2;48;85;126mj\033[38;2;52;84;124mj\033[38;2;55;82;122mj\033[38;2;55;82;121mj\033[38;2;57;81;120mj\033[38;2;58;79;117mf\033[38;2;56;78;117mff\033[38;2;55;76;114mf\033[38;2;45;67;100m?\033[38;2;46;65;95m?\033[38;2;54;76;111mt\033[38;2;54;78;111mf\033[38;2;57;80;112mf\033[38;2;39;54;77m+\033[38;2;28;45;72mi\033[38;2;58;75;104mt\033[38;2;102;107;117mv\033[38;2;182;167;148mZ\033[38;2;237;217;179mo\033[38;2;246;231;195mM\033[38;2;248;230;195mM\033[38;2;247;228;192mM\033[38;2;248;229;193mM\033[38;2;251;232;199mW\033[38;2;125;126;128mY\033[38;2;94;88;90mr\033[38;2;210;188;155mp\033[38;2;83;90;105mr\033[38;2;49;69;101m1\033[38;2;46;64;90m-\033[38;2;29;39;59m!\033[38;2;30;40;58m!\033[38;2;27;37;55ml\033[38;2;28;37;55ml\033[38;2;25;30;50mI\033[38;2;25;33;50ml\033[38;2;27;36;53ml\033[38;2;26;35;52mll\033[38;2;24;32;49mI\033[38;2;24;33;51ml\033[38;2;37;55;73m+\033[38;2;39;59;78m+\033[38;2;39;56;73m+\033[38;2;177;180;182mq\033[38;2;255;255;255m$\033[0m                   \033[0m");
  $display("\033[0m    \033[38;2;255;0;0mff\033[38;2;255;19;19mx\033[38;2;255;27;27mn\033[38;2;255;0;0mfff\033[0m      \033[38;2;255;0;0mf\033[38;2;255;223;207mW\033[38;2;255;255;255m$\033[38;2;168;183;196mp\033[38;2;69;94;129mx\033[38;2;105;125;154mY\033[38;2;180;190;204mb\033[38;2;88;110;143mc\033[38;2;56;82;124mj\033[38;2;60;86;127mr\033[38;2;58;84;125mj\033[38;2;59;85;125mj\033[38;2;54;80;117mf\033[38;2;55;79;118mf\033[38;2;58;82;122mj\033[38;2;56;82;122mjj\033[38;2;57;82;121mjj\033[38;2;56;80;120mf\033[38;2;56;78;118mf\033[38;2;57;76;117mf\033[38;2;56;78;115mf\033[38;2;54;77;112mf\033[38;2;55;76;111mt\033[38;2;45;65;97m?\033[38;2;47;66;99m?\033[38;2;50;72;107m1\033[38;2;54;79;112mf\033[38;2;52;73;104m1\033[38;2;44;50;66m~\033[38;2;158;151;140mQ\033[38;2;214;198;171mk\033[38;2;231;211;178ma\033[38;2;209;191;163md\033[38;2;195;179;157mq\033[38;2;194;180;161mq\033[38;2;196;182;162mp\033[38;2;198;184;163mp\033[38;2;199;185;162mp\033[38;2;204;189;166md\033[38;2;186;174;155mw\033[38;2;87;91;95mr\033[38;2;159;147;126mL\033[38;2;183;176;157mw\033[38;2;53;67;94m?\033[38;2;48;65;87m-\033[38;2;29;38;55ml\033[38;2;29;37;55mll\033[38;2;24;33;50mI\033[38;2;45;47;53mi\033[38;2;52;52;57m~\033[38;2;24;33;51ml\033[38;2;26;37;54ml\033[38;2;27;36;53ml\033[38;2;24;33;50mI\033[38;2;22;29;48mI\033[38;2;31;45;64mi\033[38;2;40;59;74m+\033[38;2;42;62;79m_\033[38;2;50;68;84m-\033[38;2;178;183;189mp\033[38;2;255;255;255m$$\033[0m                 \033[0m");
  $display("\033[0m      \033[38;2;255;0;0mfff\033[0m        \033[38;2;255;255;255m$\033[38;2;247;248;248mB\033[38;2;134;149;171mQ\033[38;2;77;101;137mu\033[38;2;168;180;196mp\033[38;2;255;255;255m$\033[38;2;157;171;188mw\033[38;2;56;81;120mf\033[38;2;61;84;125mr\033[38;2;58;84;124mjj\033[38;2;56;81;117mf\033[38;2;55;81;117mf\033[38;2;57;83;123mj\033[38;2;56;82;122mjj\033[38;2;56;81;120mf\033[38;2;53;76;114mf\033[38;2;57;80;117mf\033[38;2;56;78;117mf\033[38;2;56;75;116mf\033[38;2;58;75;117mf\033[38;2;58;77;116mf\033[38;2;53;73;107mt\033[38;2;52;75;107mt\033[38;2;53;76;110mt\033[38;2;70;81;105mf\033[38;2;82;92;107mr\033[38;2;49;70;101m1\033[38;2;65;79;102mf\033[38;2;103;98;90mx\033[38;2;252;234;195mW\033[38;2;253;232;192mW\033[38;2;247;227;189mM\033[38;2;246;226;189m#\033[38;2;241;222;187m#\033[38;2;233;214;182mo\033[38;2;225;207;178ma\033[38;2;217;202;173mk\033[38;2;213;197;169mb\033[38;2;217;200;174mk\033[38;2;233;216;186mo\033[38;2;223;212;181ma\033[38;2;136;130;114mY\033[38;2;191;180;157mq\033[38;2;109;111;118mv\033[38;2;39;53;77m+\033[38;2;30;39;57m!\033[38;2;29;37;56ml\033[38;2;28;36;55ml\033[38;2;30;37;51ml\033[38;2;62;57;50m+\033[38;2;118;103;85mn\033[38;2;23;28;44m;\033[38;2;27;35;53ml\033[38;2;27;34;53ml\033[38;2;25;33;51ml\033[38;2;24;29;48mI\033[38;2;27;38;55ml\033[38;2;39;58;72m+\033[38;2;44;63;77m_\033[38;2;39;61;72m+\033[38;2;54;70;89m?\033[38;2;126;136;152mJ\033[38;2;167;174;184mw\033[38;2;199;204;209ma\033[38;2;216;218;223m#\033[38;2;214;217;222m#\033[38;2;202;206;212ma\033[38;2;241;242;244m%%\033[38;2;255;255;255m$\033[0m           \033[0m");
  $display("\033[0m                \033[38;2;255;255;255m$\033[38;2;238;239;240m%%\033[38;2;109;128;155mY\033[38;2;106;127;157mY\033[38;2;214;220;229mM\033[38;2;255;255;255m$\033[38;2;181;190;206mb\033[38;2;61;85;124mr\033[38;2;58;83;123mj\033[38;2;58;84;124mj\033[38;2;57;84;124mj\033[38;2;55;82;120mf\033[38;2;55;80;115mf\033[38;2;58;83;122mj\033[38;2;57;82;122mj\033[38;2;56;82;122mj\033[38;2;56;82;121mj\033[38;2;52;76;112mt\033[38;2;53;75;108mt\033[38;2;56;78;116mf\033[38;2;57;76;118mf\033[38;2;58;75;118mf\033[38;2;57;77;115mf\033[38;2;56;78;113mf\033[38;2;50;72;106m1\033[38;2;54;77;109mt\033[38;2;49;71;102m1\033[38;2;156;151;143mQ\033[38;2;243;226;192m#\033[38;2;190;176;158mw\033[38;2;181;171;153mm\033[38;2;199;183;157mq\033[38;2;223;206;174mh\033[38;2;227;209;176ma\033[38;2;231;212;179mo\033[38;2;235;215;183mo\033[38;2;237;217;185m*\033[38;2;236;217;184m*\033[38;2;232;215;183mo\033[38;2;234;218;184m*\033[38;2;244;226;193mM\033[38;2;246;226;193mM\033[38;2;246;224;189m#\033[38;2;247;226;190mM\033[38;2;243;225;190m#\033[38;2;222;206;177mh\033[38;2;169;159;144m0\033[38;2;42;47;61m~\033[38;2;27;34;49ml\033[38;2;37;43;55mi\033[38;2;27;30;43mI\033[38;2;92;82;78mf\033[38;2;93;80;63mt\033[38;2;158;137;105mU\033[38;2;43;42;48m!\033[38;2;26;33;50ml\033[38;2;26;37;54ml\033[38;2;25;33;51ml\033[38;2;25;29;47mI\033[38;2;25;35;52ml\033[38;2;34;54;68m~\033[38;2;38;60;76m+\033[38;2;38;60;78m+\033[38;2;79;90;100mj\033[38;2;210;213;215m*\033[38;2;145;154;166m0\033[38;2;127;138;153mJ\033[38;2;141;151;165mQ\033[38;2;152;160;172mO\033[38;2;175;181;190mp\033[38;2;237;239;240m8\033[38;2;255;255;255m$\033[0m           \033[0m");
  $display("\033[0m               \033[38;2;255;255;255m$\033[38;2;237;238;238m8\033[38;2;99;119;147mz\033[38;2;122;141;168mC\033[38;2;243;244;246mB\033[38;2;255;255;255m$\033[38;2;214;217;226m#\033[38;2;76;100;138mu\033[38;2;57;80;123mj\033[38;2;57;84;124mj\033[38;2;56;86;124mj\033[38;2;56;82;121mj\033[38;2;53;78;116mf\033[38;2;57;83;122mj\033[38;2;56;82;122mj\033[38;2;57;82;122mjj\033[38;2;57;81;118mf\033[38;2;50;73;106m1\033[38;2;57;78;114mf\033[38;2;56;76;117mf\033[38;2;56;75;117mff\033[38;2;53;75;113mt\033[38;2;54;77;109mt\033[38;2;52;74;109mt\033[38;2;52;75;110mt\033[38;2;51;70;97m1\033[38;2;198;186;165mp\033[38;2;252;232;195mW\033[38;2;253;231;194mW\033[38;2;245;225;189m#\033[38;2;157;140;119mJ\033[38;2;126;112;100mv\033[38;2;126;118;107mz\033[38;2;132;127;117mX\033[38;2;165;158;147m0\033[38;2;129;121;111mz\033[38;2;118;109;97mv\033[38;2;112;100;86mn\033[38;2;150;134;118mU\033[38;2;240;223;195m#\033[38;2;242;225;195m#\033[38;2;242;224;191m###\033[38;2;246;227;194mM\033[38;2;237;218;184m*\033[38;2;187;166;134mZ\033[38;2;148;129;102mY\033[38;2;160;139;109mJ\033[38;2;148;124;96mX\033[38;2;122;103;84mn\033[38;2;116;98;78mx\033[38;2;166;143;107mJ\033[38;2;66;62;57m_\033[38;2;22;30;47mI\033[38;2;28;36;52ml\033[38;2;25;30;47mI\033[38;2;27;31;48mI\033[38;2;25;34;50ml\033[38;2;31;46;60mi\033[38;2;37;56;71m+\033[38;2;42;63;80m_\033[38;2;35;52;70m~\033[38;2;172;174;175mw\033[38;2;255;255;255m$$$$$\033[0m             \033[0m");
  $display("\033[0m              \033[38;2;255;255;255m$\033[38;2;241;241;241m%%\033[38;2;102;120;146mX\033[38;2;118;137;165mC\033[38;2;249;251;251m@\033[0m \033[38;2;255;255;255m$\033[38;2;138;153;177m0\033[38;2;49;75;116mt\033[38;2;60;84;125mj\033[38;2;57;84;124mj\033[38;2;56;85;122mj\033[38;2;52;77;114mf\033[38;2;57;84;122mj\033[38;2;56;84;123mj\033[38;2;56;82;122mj\033[38;2;57;82;122mjj\033[38;2;53;77;113mf\033[38;2;51;74;107mt\033[38;2;56;78;116mf\033[38;2;54;76;116mf\033[38;2;54;76;112mt\033[38;2;55;76;116mf\033[38;2;49;68;101m1\033[38;2;50;72;101m1\033[38;2;53;77;111mt\033[38;2;49;73;107m1\033[38;2;54;70;101m1\033[38;2;205;191;171mb\033[38;2;250;229;194mM\033[38;2;244;225;190m#\033[38;2;244;225;188m#\033[38;2;247;227;189mM\033[38;2;243;231;197mM\033[38;2;236;235;220m&\033[38;2;231;234;220mW\033[38;2;230;232;217mW\033[38;2;229;230;220mW\033[38;2;228;225;206m#\033[38;2;232;215;184mo\033[38;2;231;215;182mo\033[38;2;240;224;194m#\033[38;2;242;225;197mM\033[38;2;241;224;195m#\033[38;2;241;224;194m#\033[38;2;239;224;194m#\033[38;2;242;223;191m#\033[38;2;243;225;191m#\033[38;2;239;221;185m*\033[38;2;230;212;177ma\033[38;2;234;217;182mo\033[38;2;187;164;124mO\033[38;2;167;142;107mJ\033[38;2;170;145;112mC\033[38;2;175;148;110mL\033[38;2;74;65;60m-\033[38;2;24;28;46mI\033[38;2;30;32;49ml\033[38;2;24;30;46mI\033[38;2;24;34;50ml\033[38;2;23;33;50mI\033[38;2;26;40;56ml\033[38;2;31;50;64mi\033[38;2;44;63;79m_\033[38;2;39;58;78m+\033[38;2;89;96;107mx\033[38;2;247;245;243mB\033[0m                 \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;255;255;252m$\033[38;2;125;141;164mC\033[38;2;86;109;143mv\033[38;2;234;237;241m8\033[38;2;255;255;255m$\033[0m \033[38;2;244;244;247mB\033[38;2;94;115;146mz\033[38;2;55;81;120mf\033[38;2;59;84;124mj\033[38;2;59;85;124mj\033[38;2;54;80;114mf\033[38;2;55;80;118mf\033[38;2;57;85;125mj\033[38;2;55;83;122mj\033[38;2;56;82;122mj\033[38;2;57;82;122mj\033[38;2;56;81;121mj\033[38;2;49;73;109mt\033[38;2;54;77;112mf\033[38;2;54;77;114mf\033[38;2;54;76;113mf\033[38;2;54;76;111mt\033[38;2;55;77;114mf\033[38;2;44;61;88m-\033[38;2;45;63;91m-\033[38;2;55;80;112mf\033[38;2;49;73;106m1\033[38;2;39;60;97m-\033[38;2;161;156;149m0\033[38;2;253;233;198mW\033[38;2;244;226;191m##\033[38;2;244;225;189m#\033[38;2;238;228;199mM\033[38;2;232;232;220mW\033[38;2;230;230;218mW\033[38;2;231;231;219mW\033[38;2;231;233;220mW\033[38;2;238;230;207mW\033[38;2;242;225;190m#\033[38;2;241;225;192m#\033[38;2;241;224;194m####\033[38;2;241;224;195m#\033[38;2;240;223;191m#\033[38;2;244;225;191m#\033[38;2;232;215;185mo\033[38;2;120;106;93mu\033[38;2;130;121;105mz\033[38;2;156;141;116mJ\033[38;2;152;128;98mY\033[38;2;171;146;111mC\033[38;2;177;147;110mL\033[38;2;99;85;74mj\033[38;2;28;30;46mI\033[38;2;26;30;48mI\033[38;2;28;33;49ml\033[38;2;26;34;51ml\033[38;2;25;33;50ml\033[38;2;25;35;51ml\033[38;2;29;45;61mi\033[38;2;43;62;80m_\033[38;2;41;62;81m_\033[38;2;40;57;75m+\033[38;2;198;198;198mh\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;182;189;199mb\033[38;2;58;83;121mj\033[38;2;200;208;219mo\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;220;222;230mM\033[38;2;68;90;128mx\033[38;2;58;84;122mj\033[38;2;60;86;123mj\033[38;2;58;83;120mj\033[38;2;54;77;114mf\033[38;2;58;84;123mj\033[38;2;56;84;123mj\033[38;2;55;83;122mj\033[38;2;56;82;120mjj\033[38;2;55;81;118mf\033[38;2;48;72;106m1\033[38;2;55;76;114mf\033[38;2;55;75;114mf\033[38;2;55;77;114mf\033[38;2;54;77;113mf\033[38;2;55;78;113mf\033[38;2;42;59;85m_\033[38;2;37;50;72m~\033[38;2;55;79;111mf\033[38;2;56;76;104mt\033[38;2;125;131;137mU\033[38;2;83;91;104mr\033[38;2;223;209;184ma\033[38;2;249;232;198mW\033[38;2;242;226;192m#\033[38;2;242;225;189m#\033[38;2;236;230;204mM\033[38;2;232;232;220mW\033[38;2;232;232;219mW\033[38;2;231;233;220mW\033[38;2;232;233;218mW\033[38;2;239;226;198mM\033[38;2;241;224;194m##\033[38;2;240;223;193m#\033[38;2;240;223;192m#\033[38;2;240;223;191m#\033[38;2;241;224;192m#\033[38;2;240;224;192m#\033[38;2;241;225;194m#\033[38;2;240;226;194m#\033[38;2;242;225;189m#\033[38;2;237;217;182m*\033[38;2;202;189;162mp\033[38;2;137;136;120mU\033[38;2;76;72;64m?\033[38;2;113;98;79mx\033[38;2;168;145;106mJ\033[38;2;92;84;72mf\033[38;2;28;31;45mI\033[38;2;30;33;51ml\033[38;2;32;35;52ml\033[38;2;29;31;49ml\033[38;2;24;29;46mI\033[38;2;25;30;46mI\033[38;2;29;42;57m!\033[38;2;41;59;80m_\033[38;2;36;56;76m+\033[38;2;32;52;73m~\033[38;2;137;140;145mC\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$\033[38;2;248;248;247mB\033[38;2;90;110;138mv\033[38;2;92;115;148mz\033[38;2;250;250;251m@\033[0m  \033[38;2;255;255;255m$\033[38;2;179;186;200md\033[38;2;53;78;118mf\033[38;2;59;86;123mj\033[38;2;59;86;122mj\033[38;2;54;77;116mf\033[38;2;58;80;120mj\033[38;2;57;84;124mj\033[38;2;54;83;122mj\033[38;2;55;83;122mj\033[38;2;55;82;120mff\033[38;2;53;78;114mf\033[38;2;49;71;105m1\033[38;2;56;75;117mf\033[38;2;56;74;115mf\033[38;2;55;75;114mf\033[38;2;53;76;110mt\033[38;2;53;78;111mt\033[38;2;43;61;89m-\033[38;2;30;40;58m!\033[38;2;50;67;102m1\033[38;2;65;78;102mf\033[38;2;231;216;188mo\033[38;2;194;182;162mq\033[38;2;133;128;122mY\033[38;2;209;195;169mb\033[38;2;238;223;190m#\033[38;2;240;224;188m#\033[38;2;235;232;209mW\033[38;2;231;233;220mW\033[38;2;231;232;220mW\033[38;2;231;234;218mW\033[38;2;234;231;215mW\033[38;2;241;225;193m#\033[38;2;242;224;192m#\033[38;2;242;224;195m#\033[38;2;241;224;195m#\033[38;2;240;224;193m#\033[38;2;240;224;192m#\033[38;2;240;224;191m##\033[38;2;241;224;194m#\033[38;2;239;221;188m#\033[38;2;241;222;189m#\033[38;2;244;225;187m#\033[38;2;244;229;198mM\033[38;2;198;196;175mb\033[38;2;169;167;146mO\033[38;2;164;149;119mL\033[38;2;105;91;76mr\033[38;2;22;30;46mI\033[38;2;29;35;52ml\033[38;2;32;34;52ml\033[38;2;30;33;50ml\033[38;2;26;29;46mI\033[38;2;25;28;45mI\033[38;2;28;31;48mI\033[38;2;29;40;55m!\033[38;2;39;58;79m+\033[38;2;36;56;73m+\033[38;2;30;50;71m~\033[38;2;114;121;131mX\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$\033[38;2;238;238;239m8\033[38;2;76;98;130mn\033[38;2;75;100;135mn\033[38;2;231;233;238m8\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;141;152;174m0\033[38;2;51;76;115mt\033[38;2;58;85;122mj\033[38;2;57;81;119mf\033[38;2;52;77;116mf\033[38;2;56;83;123mj\033[38;2;55;83;122mjj\033[38;2;55;82;122mj\033[38;2;54;81;121mf\033[38;2;52;81;120mf\033[38;2;47;70;102m1\033[38;2;51;69;103m1\033[38;2;57;74;117mf\033[38;2;56;73;116mf\033[38;2;56;73;115mf\033[38;2;54;74;111mt\033[38;2;52;76;111mt\033[38;2;50;68;101m1\033[38;2;29;39;60m!\033[38;2;37;52;78m+\033[38;2;66;77;96mt\033[38;2;220;203;176mh\033[38;2;255;235;198mW\033[38;2;235;215;185mo\033[38;2;202;186;162mp\033[38;2;216;202;172mk\033[38;2;230;214;182mo\033[38;2;233;231;213mW\033[38;2;231;234;221mW\033[38;2;230;232;221mW\033[38;2;230;233;220mW\033[38;2;236;229;210mW\033[38;2;240;224;189m#\033[38;2;241;224;192m#\033[38;2;241;224;195m#\033[38;2;240;223;195m#\033[38;2;240;223;193m##\033[38;2;240;223;191m#\033[38;2;239;223;190m#\033[38;2;240;223;190m#\033[38;2;242;223;190m##\033[38;2;239;222;188m#\033[38;2;237;228;207mM\033[38;2;204;203;188mh\033[38;2;171;162;137m0\033[38;2;163;143;111mJ\033[38;2;48;46;52mi\033[38;2;28;33;51ml\033[38;2;32;35;54ml\033[38;2;29;33;51ml\033[38;2;23;30;46mI\033[38;2;23;29;46mI\033[38;2;24;32;49mI\033[38;2;25;32;49mI\033[38;2;26;39;53ml\033[38;2;40;60;76m+\033[38;2;39;58;75m+\033[38;2;34;54;68m~\033[38;2;173;176;178mw\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;148;161;178mZ\033[38;2;42;70;111m1\033[38;2;133;150;173mQ\033[38;2;255;255;255m$$$\033[38;2;165;175;192mq\033[38;2;50;76;113mt\033[38;2;59;83;120mj\033[38;2;54;77;114mf\033[38;2;55;81;120mf\033[38;2;54;83;122mj\033[38;2;55;82;121mj\033[38;2;55;83;121mj\033[38;2;55;81;120mf\033[38;2;54;80;120mf\033[38;2;52;81;118mf\033[38;2;40;57;82m_\033[38;2;50;71;105m1\033[38;2;56;74;116mf\033[38;2;56;73;116mf\033[38;2;56;73;115mf\033[38;2;54;74;110mt\033[38;2;53;76;109mt\033[38;2;54;74;108mt\033[38;2;36;47;70m~\033[38;2;29;41;61m!\033[38;2;59;67;81m?\033[38;2;198;175;145mw\033[38;2;248;232;195mW\033[38;2;244;228;191mM\033[38;2;247;229;192mM\033[38;2;244;225;188m#\033[38;2;240;227;197mM\033[38;2;232;233;220mW\033[38;2;231;233;220mWW\033[38;2;231;234;219mW\033[38;2;238;228;204mM\033[38;2;241;224;189m#\033[38;2;241;225;193m#\033[38;2;243;226;196mM\033[38;2;243;227;196mM\033[38;2;241;226;192m#\033[38;2;239;223;191m#\033[38;2;242;227;194mM\033[38;2;242;226;192m#\033[38;2;239;222;189m#\033[38;2;240;222;189m#\033[38;2;240;221;187m#\033[38;2;236;222;190m#\033[38;2;235;230;216mW\033[38;2;191;189;170mp\033[38;2;173;160;126m0\033[38;2;125;110;92mv\033[38;2;27;31;48mI\033[38;2;32;34;53ml\033[38;2;30;34;53ml\033[38;2;27;34;52ml\033[38;2;24;33;49mI\033[38;2;25;34;50ml\033[38;2;26;35;52ml\033[38;2;25;33;50ml\033[38;2;27;40;55ml\033[38;2;39;60;75m+\033[38;2;34;54;75m+\033[38;2;82;94;106mr\033[38;2;250;248;247m@\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;240;240;241m%%\033[38;2;130;146;168mL\033[38;2;51;78;116mf\033[38;2;108;127;156mY\033[38;2;175;186;201md\033[38;2;207;214;223m*\033[38;2;178;187;201md\033[38;2;58;79;115mf\033[38;2;60;80;116mf\033[38;2;52;75;111mt\033[38;2;56;82;122mj\033[38;2;55;83;122mj\033[38;2;55;82;120mf\033[38;2;56;82;119mff\033[38;2;55;82;119mf\033[38;2;51;76;109mt\033[38;2;34;47;68mi\033[38;2;52;72;107mt\033[38;2;55;74;117mf\033[38;2;55;74;116mf\033[38;2;55;74;115mf\033[38;2;54;74;112mt\033[38;2;53;75;109mt\033[38;2;53;76;111mt\033[38;2;43;61;89m-\033[38;2;27;39;57m!\033[38;2;38;48;64m~\033[38;2;140;120;100mz\033[38;2;218;195;160mb\033[38;2;245;230;196mM\033[38;2;244;227;189m#\033[38;2;242;225;188m#\033[38;2;236;229;205mM\033[38;2;232;233;222mW\033[38;2;231;232;219mW\033[38;2;230;232;219mW\033[38;2;231;233;217mW\033[38;2;240;225;194m#\033[38;2;244;224;189m#\033[38;2;240;222;191m#\033[38;2;220;197;171mk\033[38;2;197;165;141mm\033[38;2;177;140;116mL\033[38;2;160;124;106mY\033[38;2;134;110;95mc\033[38;2;213;196;170mb\033[38;2;245;226;192mM\033[38;2;239;223;189m#\033[38;2;238;223;186m*\033[38;2;237;228;203mM\033[38;2;207;207;189mh\033[38;2;174;166;139mO\033[38;2;165;148;113mC\033[38;2;59;54;54m+\033[38;2;24;30;50mI\033[38;2;29;36;54ml\033[38;2;26;35;52ml\033[38;2;25;33;51ml\033[38;2;26;31;50mI\033[38;2;26;33;51ml\033[38;2;26;35;52ml\033[38;2;25;33;50ml\033[38;2;29;42;58m!\033[38;2;40;61;77m_\033[38;2;35;57;75m+\033[38;2;33;53;69m~\033[38;2;182;187;192md\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m              \033[38;2;255;255;255m$\033[38;2;255;255;253m$\033[38;2;179;186;196md\033[38;2;103;122;148mX\033[38;2;72;96;130mn\033[38;2;73;98;132mn\033[38;2;66;91;125mr\033[38;2;59;82;115mf\033[38;2;56;79;112mf\033[38;2;52;74;110mt\033[38;2;57;82;122mj\033[38;2;56;81;121mj\033[38;2;56;82;119mff\033[38;2;55;81;118mf\033[38;2;56;81;120mf\033[38;2;44;66;94m?\033[38;2;33;43;65mi\033[38;2;54;72;109mt\033[38;2;55;74;117mf\033[38;2;55;74;116mf\033[38;2;55;74;115mf\033[38;2;54;74;112mt\033[38;2;51;73;108mt\033[38;2;52;75;110mt\033[38;2;51;72;103m1\033[38;2;34;44;62mi\033[38;2;31;40;53m!\033[38;2;28;36;47ml\033[38;2;125;107;88mu\033[38;2;200;178;145mw\033[38;2;232;213;179mo\033[38;2;244;226;190m#\033[38;2;239;232;207mW\033[38;2;234;234;222m&\033[38;2;231;232;220mW\033[38;2;230;232;220mW\033[38;2;231;233;214mW\033[38;2;241;225;191m#\033[38;2;244;223;189m#\033[38;2;192;156;132mO\033[38;2;177;127;110mJ\033[38;2;183;127;113mC\033[38;2;183;126;111mC\033[38;2;177;121;105mU\033[38;2;132;85;73mx\033[38;2;165;146;125mL\033[38;2;248;229;192mM\033[38;2;243;225;189m#\033[38;2;235;220;186m*\033[38;2;202;195;174mb\033[38;2;179;174;151mm\033[38;2;169;156;129mQ\033[38;2;86;77;73mt\033[38;2;24;29;46mI\033[38;2;30;35;52ml\033[38;2;29;35;53ml\033[38;2;27;35;53ml\033[38;2;25;31;48mI\033[38;2;26;31;50mI\033[38;2;26;33;51ml\033[38;2;26;35;52ml\033[38;2;25;32;50mI\033[38;2;31;46;62mi\033[38;2;37;56;75m+\033[38;2;64;80;95mt\033[38;2;108;123;134mz\033[38;2;72;89;103mj\033[38;2;240;240;240m%%\033[38;2;255;255;255m$\033[0m               \033[0m");
  $display("\033[0m                \033[38;2;255;255;255m$\033[38;2;252;250;247m@\033[38;2;200;204;207ma\033[38;2;171;178;184mq\033[38;2;177;185;189mp\033[38;2;199;202;208ma\033[38;2;74;93;123mx\033[38;2;50;72;110mt\033[38;2;57;83;121mj\033[38;2;57;83;120mj\033[38;2;56;83;118mf\033[38;2;55;82;118mf\033[38;2;54;80;117mf\033[38;2;55;81;118mf\033[38;2;41;58;85m_\033[38;2;32;44;63mi\033[38;2;53;72;108mt\033[38;2;53;74;114mt\033[38;2;54;74;115mf\033[38;2;54;73;115mt\033[38;2;54;74;111mt\033[38;2;51;74;108mtt\033[38;2;53;74;107mt\033[38;2;37;50;73m~\033[38;2;32;39;54m!\033[38;2;21;30;48mI\033[38;2;116;102;84mn\033[38;2;182;156;119mQ\033[38;2;181;153;119mQ\033[38;2;195;171;134mZ\033[38;2;211;196;167mb\033[38;2;225;221;205m#\033[38;2;232;234;223mW\033[38;2;232;237;225m&\033[38;2;236;233;212mW\033[38;2;244;224;188m#\033[38;2;244;224;189m#\033[38;2;235;213;180mo\033[38;2;235;209;177mo\033[38;2;237;208;177mo\033[38;2;233;201;172mh\033[38;2;225;191;163mb\033[38;2;219;189;160mb\033[38;2;233;211;178mo\033[38;2;242;221;183m*\033[38;2;217;200;168mk\033[38;2;190;179;156mw\033[38;2;170;166;147mO\033[38;2;135;133;120mY\033[38;2;63;63;64m-\033[38;2;26;29;49mI\033[38;2;31;34;54ml\033[38;2;29;32;51ml\033[38;2;28;34;52ml\033[38;2;26;32;50ml\033[38;2;25;30;47mI\033[38;2;26;33;51ml\033[38;2;25;34;52ml\033[38;2;26;35;52ml\033[38;2;25;33;48mI\033[38;2;34;52;68m~\033[38;2;29;50;70mi\033[38;2;155;161;167mO\033[38;2;255;255;255m$\033[38;2;78;91;110mr\033[38;2;164;169;178mm\033[38;2;255;255;255m$\033[0m               \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;177;185;191mp\033[38;2;54;75;107mt\033[38;2;58;82;117mf\033[38;2;58;82;119mj\033[38;2;58;81;117mff\033[38;2;57;80;117mf\033[38;2;57;79;114mf\033[38;2;39;53;78m+\033[38;2;32;44;61mi\033[38;2;50;69;104m1\033[38;2;53;76;110mt\033[38;2;53;75;112mt\033[38;2;55;73;114mt\033[38;2;55;75;111mt\033[38;2;53;76;110mt\033[38;2;52;75;109mt\033[38;2;53;76;110mt\033[38;2;43;59;84m_\033[38;2;30;36;52ml\033[38;2;37;37;51m!\033[38;2;150;129;103mY\033[38;2;184;156;118mQ\033[38;2;181;154;117mQ\033[38;2;179;153;115mQ\033[38;2;178;151;115mL\033[38;2;182;156;121m0\033[38;2;192;173;144mm\033[38;2;204;197;175mb\033[38;2;224;217;193mo\033[38;2;242;225;191m#\033[38;2;251;232;193mW\033[38;2;251;230;193mM\033[38;2;246;226;190m#\033[38;2;244;225;189m#\033[38;2;247;228;191mM\033[38;2;252;232;194mW\033[38;2;249;225;189mM\033[38;2;223;197;163mk\033[38;2;183;162;132mO\033[38;2;148;142;122mJ\033[38;2;111;109;104mv\033[38;2;62;64;71m-\033[38;2;28;34;50ml\033[38;2;25;33;52ml\033[38;2;28;34;53ml\033[38;2;29;34;53ml\033[38;2;26;31;50mI\033[38;2;27;34;52ml\033[38;2;24;31;49mI\033[38;2;25;33;50ml\033[38;2;26;35;52mll\033[38;2;26;34;52ml\033[38;2;27;38;53ml\033[38;2;28;47;66mi\033[38;2;125;136;148mJ\033[38;2;255;255;255m$$\033[38;2;165;171;183mw\033[38;2;94;103;123mu\033[38;2;255;255;255m$$\033[0m              \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;227;229;230mW\033[38;2;64;86;116mj\033[38;2;50;71;102m1\033[38;2;58;80;114mf\033[38;2;57;81;114mf\033[38;2;57;79;113mf\033[38;2;56;80;115mf\033[38;2;57;79;112mf\033[38;2;40;53;76m+\033[38;2;36;42;63mi\033[38;2;48;66;100m?\033[38;2;53;76;113mt\033[38;2;54;74;113mt\033[38;2;54;74;111mt\033[38;2;54;75;110mt\033[38;2;53;75;110mt\033[38;2;53;75;109mt\033[38;2;53;76;109mt\033[38;2;48;68;98m?\033[38;2;31;37;57m!\033[38;2;42;43;57mi\033[38;2;151;147;134mL\033[38;2;164;147;121mL\033[38;2;173;148;112mL\033[38;2;180;152;115mQ\033[38;2;181;154;116mQ\033[38;2;182;153;115mQ\033[38;2;181;152;112mL\033[38;2;178;150;111mL\033[38;2;180;155;118mQ\033[38;2;158;143;118mJ\033[38;2;136;129;117mY\033[38;2;192;176;155mw\033[38;2;228;210;180ma\033[38;2;242;222;188m#\033[38;2;221;203;171mh\033[38;2;183;165;140mZ\033[38;2;133;117;102mz\033[38;2;86;78;75mt\033[38;2;55;57;63m+\033[38;2;34;42;56m!\033[38;2;23;33;48mI\033[38;2;24;34;52ml\033[38;2;28;37;55ml\033[38;2;28;37;54ml\033[38;2;26;34;52ml\033[38;2;27;34;52ml\033[38;2;24;31;49mI\033[38;2;26;33;51ml\033[38;2;24;31;49mI\033[38;2;25;34;51ml\033[38;2;25;35;52ml\033[38;2;26;34;52ml\033[38;2;24;33;51ml\033[38;2;23;40;57ml\033[38;2;108;122;134mz\033[38;2;240;242;242m%%\033[38;2;255;255;255m$$\033[38;2;216;218;223m#\033[38;2;84;95;118mn\033[38;2;245;245;247mB\033[38;2;255;255;255m$\033[0m              \033[0m");
  $display("\033[0m                \033[38;2;251;251;251m@\033[38;2;255;255;255m$$\033[0m \033[38;2;255;255;255m$$\033[38;2;150;163;182mZ\033[38;2;62;87;122mr\033[38;2;53;75;103mt\033[38;2;41;58;85m_\033[38;2;48;68;103m1\033[38;2;57;80;116mf\033[38;2;57;80;113mf\033[38;2;57;79;114mf\033[38;2;42;55;80m_\033[38;2;37;42;61mi\033[38;2;44;59;85m_\033[38;2;54;77;114mf\033[38;2;53;75;113mt\033[38;2;53;75;112mt\033[38;2;53;76;110mt\033[38;2;52;74;109mt\033[38;2;52;75;109mt\033[38;2;51;74;108mt\033[38;2;51;73;107mt\033[38;2;39;51;77m+\033[38;2;25;31;49mI\033[38;2;122;128;129mY\033[38;2;170;176;163mm\033[38;2;159;157;142mQ\033[38;2;161;146;123mC\033[38;2;171;147;113mC\033[38;2;180;151;112mL\033[38;2;181;154;114mQ\033[38;2;182;153;114mQ\033[38;2;180;152;113mL\033[38;2;103;95;88mx\033[38;2;21;28;47mI\033[38;2;34;40;57m!\033[38;2;56;62;71m-\033[38;2;71;75;82m1\033[38;2;48;53;61m+\033[38;2;30;39;52ml\033[38;2;24;35;51ml\033[38;2;25;35;53ml\033[38;2;29;37;56ml\033[38;2;30;37;55ml\033[38;2;29;38;52ml\033[38;2;29;37;55ml\033[38;2;29;38;55ml\033[38;2;26;35;52ml\033[38;2;26;34;51ml\033[38;2;27;34;52ml\033[38;2;23;30;48mI\033[38;2;26;33;51ml\033[38;2;26;35;52mll\033[38;2;26;34;52ml\033[38;2;24;32;48mI\033[38;2;20;31;49mI\033[38;2;95;108;123mv\033[38;2;241;242;242m%%\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;173;179;189mp\033[38;2;109;118;137mz\033[38;2;255;255;255m$$\033[0m              \033[0m");
  $display("\033[0m               \033[38;2;255;255;255m$$\033[38;2;241;244;248mB\033[38;2;202;209;219mo\033[38;2;191;200;211mh\033[38;2;184;192;206mk\033[38;2;152;167;189mm\033[38;2;142;157;178mO\033[38;2;174;184;199md\033[38;2;56;81;116mf\033[38;2;110;122;133mz\033[38;2;105;113;121mc\033[38;2;46;62;88m-\033[38;2;54;76;107mt\033[38;2;57;82;115mf\033[38;2;47;60;87m-\033[38;2;39;45;62mi\033[38;2;39;53;72m+\033[38;2;54;76;112mt\033[38;2;53;76;112mt\033[38;2;53;77;111mt\033[38;2;53;76;110mt\033[38;2;53;76;109mtt\033[38;2;51;74;108mt\033[38;2;51;74;109mt\033[38;2;47;67;98m?\033[38;2;27;36;57ml\033[38;2;54;59;70m_\033[38;2;161;165;155mO\033[38;2;171;175;165mm\033[38;2;166;169;161mZ\033[38;2;160;159;147m0\033[38;2;160;147;125mL\033[38;2;169;146;112mC\033[38;2;179;150;109mL\033[38;2;164;141;109mJ\033[38;2;157;160;150m0\033[38;2;98;102;102mn\033[38;2;27;36;52ml\033[38;2;31;40;59m!\033[38;2;30;40;58m!\033[38;2;31;41;59m!\033[38;2;31;39;57m!\033[38;2;30;37;55ml\033[38;2;29;36;54ml\033[38;2;32;38;57m!\033[38;2;30;37;54ml\033[38;2;29;38;52ml\033[38;2;29;37;56ml\033[38;2;28;37;55ml\033[38;2;25;33;52ml\033[38;2;25;32;51ml\033[38;2;23;30;49mI\033[38;2;23;31;49mI\033[38;2;26;34;52ml\033[38;2;26;35;52mll\033[38;2;25;33;50ml\033[38;2;22;34;50mI\033[38;2;47;62;81m-\033[38;2;213;214;219m*\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;223;224;228mW\033[38;2;82;93;115mx\033[38;2;212;216;222m#\033[38;2;255;255;255m$\033[0m               \033[0m");
  $display("\033[0m                \033[38;2;255;255;255m$\033[38;2;246;246;250mB\033[38;2;218;222;231mM\033[38;2;200;207;217mo\033[38;2;194;203;214ma\033[38;2;210;216;222m#\033[38;2;255;255;255m$\033[38;2;116;135;163mJ\033[38;2;144;158;175mO\033[38;2;255;255;253m$\033[38;2;255;255;255m$\033[38;2;125;133;140mU\033[38;2;31;44;67mi\033[38;2;45;63;93m-\033[38;2;53;68;98m1\033[38;2;40;46;66m~\033[38;2;37;47;62mi\033[38;2;52;69;100m1\033[38;2;54;77;115mf\033[38;2;53;76;111mt\033[38;2;53;76;110mt\033[38;2;54;77;111mt\033[38;2;53;76;110mt\033[38;2;50;73;107m1\033[38;2;51;72;107m1\033[38;2;52;75;108mt\033[38;2;40;56;84m_\033[38;2;24;32;56ml\033[38;2;76;80;88mf\033[38;2;164;169;156mZ\033[38;2;172;176;160mm\033[38;2;168;172;159mZ\033[38;2;168;171;160mZ\033[38;2;159;159;149m0\033[38;2;156;148;130mL\033[38;2;150;145;128mC\033[38;2;149;153;143mL\033[38;2;167;170;159mZ\033[38;2;81;88;90mj\033[38;2;31;38;55m!\033[38;2;29;37;55ml\033[38;2;33;41;59m!\033[38;2;32;39;58m!\033[38;2;29;36;55ml\033[38;2;29;37;55mll\033[38;2;29;38;54mll\033[38;2;28;38;55ml\033[38;2;28;37;56ml\033[38;2;24;32;51mI\033[38;2;22;29;48mI\033[38;2;24;32;51mI\033[38;2;25;34;51ml\033[38;2;26;35;52ml\033[38;2;25;34;51ml\033[38;2;24;34;51ml\033[38;2;28;40;58m!\033[38;2;27;45;66mi\033[38;2;115;122;130mX\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;199;203;211ma\033[38;2;94;105;126mv\033[38;2;165;170;182mw\033[38;2;255;255;255m$$\033[0m               \033[0m");
  $display("\033[0m                      \033[38;2;255;255;255m$\033[38;2;129;147;173mQ\033[38;2;181;191;206mb\033[38;2;255;255;255m$\033[38;2;253;252;250m@\033[38;2;146;154;159m0\033[38;2;90;103;117mn\033[38;2;72;79;92mf\033[38;2;37;48;70m~\033[38;2;43;51;73m+\033[38;2;42;48;66m~\033[38;2;45;55;82m_\033[38;2;55;76;114mf\033[38;2;52;76;112mt\033[38;2;54;77;111mtt\033[38;2;53;77;111mt\033[38;2;52;75;107mt\033[38;2;45;64;93m-\033[38;2;47;63;92m-\033[38;2;52;72;106m1\033[38;2;38;52;77m+\033[38;2;26;33;53ml\033[38;2;64;70;79m?\033[38;2;149;152;143mL\033[38;2;172;174;160mm\033[38;2;168;170;156mZ\033[38;2;155;158;149m0\033[38;2;149;155;149mQ\033[38;2;145;152;144mL\033[38;2;151;157;146mQ\033[38;2;163;166;155mO\033[38;2;121;125;118mz\033[38;2;107;115;115mv\033[38;2;65;72;78m?\033[38;2;36;41;56m!\033[38;2;26;33;51ml\033[38;2;26;33;53ml\033[38;2;30;39;57m!\033[38;2;29;38;55mll\033[38;2;29;37;55ml\033[38;2;27;36;53ml\033[38;2;23;32;50mI\033[38;2;23;30;49mI\033[38;2;26;32;50ml\033[38;2;26;35;52ml\033[38;2;25;35;52ml\033[38;2;26;35;52ml\033[38;2;25;34;52ml\033[38;2;26;35;54ml\033[38;2;27;41;56m!\033[38;2;28;48;63mi\033[38;2;145;147;149mL\033[38;2;252;252;253m$\033[38;2;183;187;196md\033[38;2;148;155;169m0\033[38;2;127;136;154mJ\033[38;2;197;201;207mh\033[38;2;255;255;255m$\033[0m                 \033[0m");
  $display("\033[0m                      \033[38;2;255;255;255m$\033[38;2;238;242;245m%%\033[38;2;208;214;221m*\033[38;2;245;244;238m%%\033[38;2;224;223;212m#\033[38;2;210;210;198ma\033[38;2;244;242;229m8\033[38;2;224;223;211m#\033[38;2;90;93;100mr\033[38;2;38;44;67mi\033[38;2;45;52;75m+\033[38;2;42;49;66m~\033[38;2;49;65;91m?\033[38;2;54;79;113mf\033[38;2;54;77;110mt\033[38;2;50;73;108mt\033[38;2;49;73;107m1\033[38;2;53;76;110mt\033[38;2;50;74;106m1\033[38;2;39;54;78m+\033[38;2;39;50;74m+\033[38;2;48;65;94m?\033[38;2;37;49;71m~\033[38;2;29;37;55ml\033[38;2;59;69;81m?\033[38;2;108;117;121mc\033[38;2;138;141;134mJ\033[38;2;165;169;158mZ\033[38;2;156;160;149m0\033[38;2;157;161;150m0\033[38;2;157;162;153m0\033[38;2;133;144;143mC\033[38;2;77;94;112mr\033[38;2;72;99;123mx\033[38;2;109;126;131mX\033[38;2;145;148;142mL\033[38;2;110;114;112mv\033[38;2;53;59;69m_\033[38;2;27;35;54ml\033[38;2;31;40;57m!\033[38;2;30;38;56m!\033[38;2;28;35;53ml\033[38;2;24;31;49mI\033[38;2;25;32;50mI\033[38;2;26;35;52ml\033[38;2;25;35;52mll\033[38;2;26;35;52mlll\033[38;2;24;33;50mI\033[38;2;22;36;51ml\033[38;2;25;47;61m!\033[38;2;105;106;110mu\033[38;2;251;251;250m@\033[38;2;191;194;203mk\033[38;2;198;202;210ma\033[38;2;255;255;255m$$\033[0m                  \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;253;253;250m$\033[38;2;247;245;236m%%\033[38;2;245;243;231m%%\033[38;2;238;237;225m&\033[38;2;239;239;227m8\033[38;2;241;241;228m8\033[38;2;239;238;226m8\033[38;2;244;243;229m8\033[38;2;224;225;215mM\033[38;2;80;84;93mf\033[38;2;42;49;67m~\033[38;2;43;51;70m+\033[38;2;41;49;67m~\033[38;2;48;67;95m?\033[38;2;49;73;107m1\033[38;2;90;103;124mu\033[38;2;80;93;116mx\033[38;2;44;65;100m?\033[38;2;51;74;106mt\033[38;2;53;72;103m1\033[38;2;38;51;71m~\033[38;2;33;43;63mi\033[38;2;43;56;82m_\033[38;2;36;46;67mi\033[38;2;31;40;58m!\033[38;2;55;76;99m1\033[38;2;75;100;122mn\033[38;2;99;118;129mc\033[38;2;118;130;131mY\033[38;2;129;139;139mJ\033[38;2;92;108;119mu\033[38;2;69;95;119mr\033[38;2;73;100;126mn\033[38;2;72;101;126mn\033[38;2;78;100;117mx\033[38;2;159;164;157mO\033[38;2;173;178;164mw\033[38;2;136;141;133mJ\033[38;2;30;39;50ml\033[38;2;30;39;56m!\033[38;2;29;36;54ml\033[38;2;27;34;52ml\033[38;2;27;37;54ml\033[38;2;26;38;54mlll\033[38;2;26;37;53ml\033[38;2;26;35;52ml\033[38;2;27;36;53mll\033[38;2;21;30;47mI\033[38;2;82;88;97mj\033[38;2;89;103;116mn\033[38;2;32;49;65mi\033[38;2;140;153;162mQ\033[38;2;224;229;231mW\033[38;2;212;217;222m#\033[38;2;187;195;201mk\033[38;2;225;229;232mW\033[38;2;255;255;255m$\033[0m                 \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;251;251;249m@\033[38;2;248;248;236mB\033[38;2;237;237;224m&\033[38;2;239;239;227m8\033[38;2;238;238;227m8\033[38;2;237;237;225m&\033[38;2;236;237;223m&\033[38;2;237;238;224m&\033[38;2;238;239;225m8\033[38;2;247;248;232m%%\033[38;2;179;180;175mq\033[38;2;40;44;62mi\033[38;2;50;54;72m+\033[38;2;42;48;65m~\033[38;2;40;51;69m~\033[38;2;40;60;88m_\033[38;2;72;89;112mr\033[38;2;202;205;201mh\033[38;2;96;106;122mv\033[38;2;43;63;94m-\033[38;2;50;69;104m1\033[38;2;50;72;100m1\033[38;2;33;47;67mi\033[38;2;32;42;61mi\033[38;2;42;50;71m+\033[38;2;34;40;58m!\033[38;2;37;47;66m~\033[38;2;70;93;118mr\033[38;2;69;98;124mx\033[38;2;66;92;120mr\033[38;2;60;85;110mf\033[38;2;67;91;115mr\033[38;2;68;90;112mr\033[38;2;74;99;122mx\033[38;2;71;99;124mx\033[38;2;66;93;120mr\033[38;2;107;116;115mv\033[38;2;164;165;150mO\033[38;2;166;168;158mZ\033[38;2;61;68;72m-\033[38;2;25;33;50ml\033[38;2;30;37;55mll\033[38;2;29;38;55mll\033[38;2;27;37;54ml\033[38;2;26;38;54mllll\033[38;2;26;36;54ml\033[38;2;15;23;43m;\033[38;2;121;125;129mX\033[38;2;248;247;247mB\033[38;2;157;165;173mZ\033[38;2;105;123;137mz\033[38;2;123;139;152mJ\033[38;2;137;151;162mQ\033[38;2;145;157;166m0\033[38;2;217;221;225mM\033[38;2;255;255;255m$\033[0m                 \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;252;250;250m@\033[38;2;241;239;227m8\033[38;2;225;225;209m#\033[38;2;228;226;213mM\033[38;2;227;226;215mM\033[38;2;235;235;223m&\033[38;2;237;237;225m&\033[38;2;237;238;224m&\033[38;2;234;235;220mW\033[38;2;233;233;218mW\033[38;2;242;242;230m8\033[38;2;159;159;157mO\033[38;2;55;57;69m_\033[38;2;183;183;181mp\033[38;2;86;92;99mr\033[38;2;26;35;52ml\033[38;2;70;76;88mt\033[38;2;114;125;141mY\033[38;2;124;131;141mU\033[38;2;229;230;218mW\033[38;2;163;167;165mZ\033[38;2;75;85;108mj\033[38;2;44;63;95m-\033[38;2;43;60;88m-\033[38;2;34;43;62mi\033[38;2;35;43;61mi\033[38;2;36;43;62mi\033[38;2;34;38;55m!\033[38;2;49;62;83m-\033[38;2;70;95;120mx\033[38;2;87;105;121mu\033[38;2;119;130;132mY\033[38;2;135;142;137mJ\033[38;2;134;140;132mJ\033[38;2;134;143;138mJ\033[38;2;106;106;83mx\033[38;2;109;105;72mx\033[38;2;123;108;57mx\033[38;2;141;129;84mz\033[38;2;163;164;151mO\033[38;2;133;135;128mU\033[38;2;42;44;57mi\033[38;2;33;36;56m!\033[38;2;31;38;56m!\033[38;2;28;38;53ml\033[38;2;27;38;53ml\033[38;2;29;37;54ml\033[38;2;29;36;54ml\033[38;2;29;37;53ml\033[38;2;27;35;52ml\033[38;2;22;31;48mI\033[38;2;29;36;47ml\033[38;2;27;31;41mI\033[38;2;83;88;90mj\033[38;2;255;255;255m$$$$$$\033[0m                   \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;248;247;242mB\033[38;2;236;236;220m&\033[38;2;237;238;220m&\033[38;2;237;238;222m&\033[38;2;233;233;216mW\033[38;2;223;221;206m#\033[38;2;234;233;220mW\033[38;2;239;240;226m8\033[38;2;234;234;221mW\033[38;2;225;226;213mM\033[38;2;212;212;201mo\033[38;2;161;161;153mO\033[38;2;209;210;198ma\033[38;2;246;246;229m%%\033[38;2;216;217;206m*\033[38;2;109;113;114mv\033[38;2;55;57;69m_\033[38;2;180;180;173mq\033[38;2;169;171;168mm\033[38;2;120;125;129mX\033[38;2;187;190;183md\033[38;2;219;220;207m*\033[38;2;162;166;166mZ\033[38;2;78;93;111mr\033[38;2;39;53;75m+\033[38;2;35;43;60mi\033[38;2;38;43;59mi\033[38;2;40;42;60mi\033[38;2;38;42;53m!\033[38;2;109;102;58mj\033[38;2;140;123;67mv\033[38;2;153;145;106mU\033[38;2;147;147;126mC\033[38;2;152;154;131mL\033[38;2;136;123;81mc\033[38;2;151;125;52mv\033[38;2;154;128;52mv\033[38;2;153;127;53mv\033[38;2;146;120;50mu\033[38;2;139;128;87mz\033[38;2;168;169;156mZ\033[38;2;98;100;100mn\033[38;2;29;30;46mI\033[38;2;37;39;55m!\033[38;2;35;37;53m!\033[38;2;32;36;52ml\033[38;2;32;35;52ml\033[38;2;31;33;51ml\033[38;2;25;28;46mI\033[38;2;34;37;50ml\033[38;2;63;67;66m-\033[38;2;75;79;55m?\033[38;2;24;30;24m,\033[38;2;107;113;106mv\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;252;252;244m@\033[38;2;236;238;222m&\033[38;2;237;238;220m&\033[38;2;236;237;219m&\033[38;2;239;239;220m&\033[38;2;235;233;217mW\033[38;2;191;190;177md\033[38;2;223;224;208m#\033[38;2;237;239;222m&\033[38;2;236;238;222m&\033[38;2;235;237;222m&\033[38;2;241;243;225m8\033[38;2;237;239;222m&\033[38;2;233;234;218mW\033[38;2;238;239;222m&\033[38;2;239;240;223m8\033[38;2;208;209;196ma\033[38;2;188;188;174mp\033[38;2;231;231;215mW\033[38;2;218;218;206m*\033[38;2;144;151;153mQ\033[38;2;109;119;127mz\033[38;2;136;140;144mC\033[38;2;136;142;145mC\033[38;2;62;72;82m1\033[38;2;35;42;59mi\033[38;2;41;45;60mi\033[38;2;41;44;60mi\033[38;2;33;36;47ml\033[38;2;161;142;82mY\033[38;2;190;164;74mC\033[38;2;157;133;51mc\033[38;2;139;116;50mn\033[38;2;138;116;49mn\033[38;2;141;115;50mn\033[38;2;142;118;53mu\033[38;2;150;126;52mv\033[38;2;150;125;51mv\033[38;2;151;125;50mv\033[38;2;146;122;46mu\033[38;2;146;134;95mX\033[38;2;129;132;125mY\033[38;2;32;35;48ml\033[38;2;36;37;53m!\033[38;2;38;39;55m!\033[38;2;33;37;52ml\033[38;2;30;33;48ml\033[38;2;39;43;54mi\033[38;2;73;79;84mt\033[38;2;125;129;129mY\033[38;2;135;139;131mJ\033[38;2;61;64;56m_\033[38;2;48;52;43mi\033[38;2;193;194;188mb\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;252;252;251m@\033[38;2;247;245;232m%%\033[38;2;236;237;219m&\033[38;2;234;237;219m&\033[38;2;234;237;218mW\033[38;2;236;238;220m&\033[38;2;233;232;216mW\033[38;2;183;183;170mq\033[38;2;189;190;176md\033[38;2;225;225;208m#\033[38;2;236;238;220m&\033[38;2;235;238;220m&\033[38;2;234;237;220m&\033[38;2;232;235;218mW\033[38;2;233;234;217mW\033[38;2;232;233;217mW\033[38;2;232;234;216mW\033[38;2;235;238;218m&\033[38;2;236;238;219m&\033[38;2;232;235;215mW\033[38;2;234;236;217mW\033[38;2;239;241;222m8\033[38;2;223;226;212m#\033[38;2;186;189;181md\033[38;2;154;157;154m0\033[38;2;103;108;110mu\033[38;2;35;42;55m!\033[38;2;42;47;62m~\033[38;2;42;44;61mi\033[38;2;32;35;47ml\033[38;2;176;156;90mC\033[38;2;239;211;104mp\033[38;2;227;200;93mw\033[38;2;195;171;81mQ\033[38;2;147;128;85mz\033[38;2;149;143;115mJ\033[38;2;136;136;116mY\033[38;2;145;144;114mU\033[38;2;146;137;95mY\033[38;2;146;132;80mz\033[38;2;134;118;68mu\033[38;2;117;106;61mr\033[38;2;144;148;128mC\033[38;2;108;113;108mv\033[38;2;41;43;53mi\033[38;2;29;33;48ml\033[38;2;31;37;52ml\033[38;2;32;36;50ml\033[38;2;61;67;72m-\033[38;2;72;79;79m1\033[38;2;86;90;91mj\033[38;2;83;87;88mj\033[38;2;90;93;86mj\033[38;2;203;203;197mh\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;250;250;247m@\033[38;2;243;242;224m8\033[38;2;235;237;219m&\033[38;2;235;237;217mW\033[38;2;235;236;217mW\033[38;2;237;237;217m&\033[38;2;233;234;215mW\033[38;2;184;187;170mp\033[38;2;206;207;189mh\033[38;2;231;229;211mM\033[38;2;222;220;202m*\033[38;2;236;236;218m&\033[38;2;235;238;221m&\033[38;2;232;235;218mW\033[38;2;232;233;215mW\033[38;2;233;234;216mWWWWW\033[38;2;234;235;216mW\033[38;2;226;227;209m#\033[38;2;214;214;197mo\033[38;2;228;226;213mM\033[38;2;219;216;205m*\033[38;2;112;113;113mv\033[38;2;31;35;51ml\033[38;2;32;40;56m!\033[38;2;57;60;66m_\033[38;2;107;100;71mr\033[38;2;213;190;96mZ\033[38;2;217;198;104mw\033[38;2;183;175;119mO\033[38;2;201;201;175mb\033[38;2;219;220;205m*\033[38;2;203;203;190mh\033[38;2;192;194;180md\033[38;2;159;164;153mO\033[38;2;143;152;147mL\033[38;2;101;116;123mc\033[38;2;73;97;116mx\033[38;2;68;90;114mr\033[38;2;109;121;121mz\033[38;2;167;169;153mZ\033[38;2;146;145;136mC\033[38;2;110;112;106mv\033[38;2;52;56;63m+\033[38;2;31;36;50ml\033[38;2;50;57;65m+\033[38;2;59;67;70m-\033[38;2;99;105;103mn\033[38;2;121;127;119mX\033[38;2;117;118;108mc\033[38;2;205;204;197mh\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;248;247;241mB\033[38;2;236;238;218m&\033[38;2;235;237;218m&\033[38;2;235;235;215mW\033[38;2;236;235;215mW\033[38;2;237;236;216mW\033[38;2;236;237;217m&\033[38;2;188;192;174mp\033[38;2;211;213;193ma\033[38;2;240;238;219m&\033[38;2;223;220;201m*\033[38;2;187;186;168mp\033[38;2;230;231;215mW\033[38;2;234;235;218mW\033[38;2;232;233;215mWW\033[38;2;233;234;216mWWWWW\033[38;2;232;233;215mW\033[38;2;213;214;195mo\033[38;2;198;197;183mb\033[38;2;166;165;156mZ\033[38;2;122;122;117mz\033[38;2;115;117;114mc\033[38;2;141;144;138mC\033[38;2;199;200;189mk\033[38;2;158;164;138m0\033[38;2;160;176;153mZ\033[38;2;130;163;169m0\033[38;2;116;161;186m0\033[38;2;126;168;191mO\033[38;2;139;174;191mm\033[38;2;145;169;177mZ\033[38;2;168;189;194mp\033[38;2;139;165;173mO\033[38;2;100;134;153mY\033[38;2;82;114;138mv\033[38;2;73;101;122mx\033[38;2;72;100;120mx\033[38;2;80;99;112mx\033[38;2;145;151;140mL\033[38;2;160;163;149m0\033[38;2;159;163;150m0\033[38;2;98;100;97mx\033[38;2;35;35;45ml\033[38;2;137;141;131mJ\033[38;2;123;127;115mz\033[38;2;124;127;117mX\033[38;2;127;130;118mX\033[38;2;136;138;124mU\033[38;2;189;189;176mp\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m                 \033[38;2;255;255;255m$\033[38;2;253;253;255m$\033[38;2;247;247;235mB\033[38;2;233;236;217mW\033[38;2;235;235;217mW\033[38;2;236;235;217mW\033[38;2;234;235;216mW\033[38;2;234;235;217mW\033[38;2;237;238;220m&\033[38;2;200;201;182mk\033[38;2;215;216;198mo\033[38;2;235;237;217mW\033[38;2;226;228;206m#\033[38;2;168;170;150mZ\033[38;2;180;181;163mw\033[38;2;225;224;206m#\033[38;2;235;235;216mW\033[38;2;233;234;215mWW\033[38;2;233;234;216mW\033[38;2;234;235;216mWW\033[38;2;233;234;215mW\033[38;2;232;233;214mW\033[38;2;234;235;216mW\033[38;2;227;229;210mM\033[38;2;223;225;207m#\033[38;2;225;227;207m#\033[38;2;231;231;212mM\033[38;2;240;241;220m&\033[38;2;238;239;217m&\033[38;2;186;200;196mk\033[38;2;121;162;184m0\033[38;2;123;170;193mZ\033[38;2;126;171;193mZ\033[38;2;124;170;192mZ\033[38;2;123;170;192mO\033[38;2;121;166;190mO\033[38;2;105;147;167mJ\033[38;2;122;162;178m0\033[38;2;124;160;173mQ\033[38;2;126;167;181mO\033[38;2;111;147;167mC\033[38;2;89;120;140mc\033[38;2;73;98;120mx\033[38;2;104;115;119mv\033[38;2;140;143;129mJ\033[38;2;109;113;104mv\033[38;2;95;97;90mr\033[38;2;99;103;95mn\033[38;2;141;148;134mC\033[38;2;149;152;132mL\033[38;2;163;165;145m0\033[38;2;162;165;145m0\033[38;2;158;162;143m0\033[38;2;161;164;145m0\033[38;2;241;241;239m%%\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                 \033[38;2;255;255;255m$\033[38;2;252;252;249m@\033[38;2;240;239;223m8\033[38;2;241;241;223m8\033[38;2;237;238;221m&\033[38;2;237;237;221m&&\033[38;2;238;239;221m&\033[38;2;240;241;224m8\033[38;2;221;222;206m#\033[38;2;227;228;213mM\033[38;2;236;238;222m&\033[38;2;232;234;217mW\033[38;2;202;204;187mk\033[38;2;198;198;183mb\033[38;2;208;206;190mh\033[38;2;236;235;220m&\033[38;2;238;237;221m&\033[38;2;236;235;218mW\033[38;2;237;237;222m&\033[38;2;238;239;223m&&\033[38;2;237;237;221m&\033[38;2;236;237;221m&\033[38;2;232;233;216mW\033[38;2;205;206;190mh\033[38;2;201;202;187mk\033[38;2;203;205;189mh\033[38;2;222;223;207m#\033[38;2;238;239;225m8\033[38;2;236;236;219m&\033[38;2;237;234;220m&\033[38;2;192;203;202mh\033[38;2;177;199;205mbb\033[38;2;177;200;204mb\033[38;2;176;198;202mb\033[38;2;177;197;200mb\033[38;2;192;199;194mk\033[38;2;214;215;199mo\033[38;2;211;210;191ma\033[38;2;203;206;187mh\033[38;2;197;204;195mh\033[38;2;188;199;198mk\033[38;2;175;184;189mp\033[38;2;166;170;168mm\033[38;2;208;205;192mh\033[38;2;214;212;201mo\033[38;2;218;215;202mo\033[38;2;221;219;207m*\033[38;2;203;204;198mh\033[38;2;206;206;198ma\033[38;2;209;208;200ma\033[38;2;210;212;204mo\033[38;2;209;210;202mo\033[38;2;203;203;193mh\033[38;2;240;240;237m%%\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$$\033[38;2;255;255;251m$\033[38;2;255;255;250m$\033[38;2;255;255;255m$$\033[38;2;255;255;250m$\033[38;2;251;251;251m@\033[38;2;255;255;255m$$$$$$$$$\033[38;2;255;255;250m$\033[38;2;255;255;255m$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$\033[0m                         \033[0m");
endtask

endmodule